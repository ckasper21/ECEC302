`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZaHwYgb52yTRF39SHhir41dSZIHw3eXv1mpXzlCdHhK9gC3JZxdmcMIvNsSMiDIVLGcOMFbLs5ST
28oJ0kNjpA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e/eI4hkg/iRsenUGwQ2qsvZlLRfgcwOL7C10MjmIb+cZ1EKUsjTgIe8RNcRZ2UwW2jTY9+lq4vkU
dgePhwBzi3NPH+Eyleufb7OuwE9Y5b4aAQP8BUN/N+gOGzMgSo/M7p9xcM7VEB0Km45ru87i9ZI4
9o1F7ABmIucQoiPGh9A=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xeM1L2cYwW/LtubztJlVEhrHvwTYzMBTwZFaaf7VzOfQtmYe4jnO/Xhw/i7H2lYhgdrl4h8o2Y43
Wi+MuGeTry0f5/h2tuyaLI8QNBkCoggTe/RG1BNnyeYoOVX8W4NyijXEMqyXKFNyeXfft8/3l02H
3Nx2yWEa7VpJNiOgKZI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OC7xB+G+HPHBWalw4945Uz2BKnHek4LJVt6ibmwPv2acgql5SFWLmVd6rfOTc467hEESlLuSV6tB
+XBJ/HIR0hTSrH/u7AY0mkO3eIy61VGLUdC4fC+8VrNwxh4DzH6sY2LW28s7uCKPi7qz37IEyuX1
JMJE8JOud4Di39rgcEnPRcSqctWv8k799QSEgGwMrjN2meWieoKjtvufPCCCQ03nY+EHUSltEjn3
7t6PSVEXld8fTI/kBkcrgTKQhtP3IbWANh2SQgLAiphKVqKXgJRMhEFh6e0NuJeKlUPXrAeFtKe2
Ah7ABemIO0FLrhInMyGoCh2C8k/DqDB58Pe+1Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aDXEHCaDjzZjsAGZqFjZvsfjuqhCRKSxRd8m3q1zfa0pi0a7lVl3lupO/ykY4c8BDIRmw6qhH9Rs
hNDbpBc8PfaN1rx65zgzYIXcaS3/lLBKmGFq3ArgyhPPzQFXXh2+2QKvxINXLwuFLInlIoGQdR5d
s/4IrZyDjcmuZxNFf9FYDxzfaYXAXWNYQYM3hzWv1dNkVXtqNYNCPNr7wx9ObGFJ6p4KAIjVtHk1
LtM7aefXpMIy0BMLGMx+LUrtGvPnBh4T3PDHMtYNb/l+64blYczpM4KK0xCSbXHZ7eWolFSOBKjq
Mjm4kZCW6JAhwdQB5sPaQPakBj6Kyb3TkiOlFQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lqiIzLLvreibRO905o7KX6gEUh+tTK5T2DYY760VdQVA+bUmv95DalWdyBW6mQT5U1xYuH4xQrDu
nCsHkOTMacPqvlAAqAty/qvqaBRO7w8MsRDBAGKJvxpr5rqWF/SEG7ACXn764dS5MyqB14r7i/Ko
F62nH0pRgvkT+DS9FWd/5Ago4AfKg7d8h/+OpFHrkjlTz62tj1TdUPwrsBXHabiP+3TehpjbEESy
whRvuvWw/fjQXJD5966itWm9jB7soL5jvI4UWMa1bE8/9ganE3akrLwKPMUd++haU4KcNCTJbtbU
IRlmgsWQF/KULMHD58CbOUjMqeU764j1r5jtTg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52672)
`protect data_block
04GCFudQxdRb+Y9/SzkNHZvdnbPv3fO6P3I3D/8zLzYJbdJDNfYdOk+pZXHB1MPy30BMFWg89GWr
pEOfBSDLb/9xOPoGXFzdMdCjEq+m9+fvQ2b3WYJQ8HHSozOfsLMJSQXFNT5JjAgyapwcpOERDTqA
TL25b8AEoqDKUjiMcAVoIupqJYRQqh8+9hH8MTkHqziOIC5yunKbvaE8Yz0NcgYL2ngBZ+SReSCW
UkhksTt5dHGMT4W98+fmAjsxLvyBC83UUXnzEpyHyK+4J9nE+8N7pO+sSpwYqf9pqahJdF/LfjLO
3V5OaPw1wNEi5HmxyXo1VOXNHKYTB5mvAMpZiIdiD4elVi2UwjPlgrDmSRDpFLBamdcIl7gStoLd
dh2Vdn9hrVR+86lsG/7u+dHgGO/1uP2TPUbJhWZ6SY53BDDQw92ararXLYALpEQpjRGZmr/W75SL
bwzQtEZOKKLtZTVojdvZS8qB/biT2B/THFXKp8t/wDKfUcV6TxMdLze21MgMn+NXVILH6lLsa6L8
Hmge5ter8GRXuQDX/PVP1llWLqS0yVb0/FwkhzyjQjQ5L9U7S9lnyh1Ou3ZaTg0HLrSGowhe4Rts
hPG0YXX4CXBYHAwviqf7EkUuiKoo5Q6njYTjeg926TZB7+7fkllAukWYEB+qqT9J6+HXyguGbcnr
OmujF1I7MD1eFUcn+LGXb6Bzqps0i3afxSB8onXkTtYcDEETHFRMBMYRk9E3IR2gRy1wAPpqcsgI
lTzx3fcUP3eeRPjEdadntitwZYPOObnbF0kAa0+1hxseamzBpzIz0T1hAYyofvWncuxSQULPU9p8
hmeEqK/u20Dr0zUKEqHgLAHey8fMdhcGp4RYLO4TSy7nOHpAqDy6KqfRyI3IKirxbTmTuJI6U2Dk
hRdeM10dsV3+j9qeGHm6T4kNWkr5T0Ghru3wvZE6E5IG19TzkaedGwdK/zmdOJL75nZuYWHmPExw
1cgbL4G9xUKKHnkylmAq4Ughq4cMn0rft8xLKf/HMgZ9ZIKr2yf6rxSHClbjTY7tWHn23i9YuSNO
2V36fBoli4RaQ23aP1TxQLoqMZzGGRf/v2XiZ8N3fRuhhGLqgdfXhpqOoAEqmsnYYHNCmh2JyGzt
V4VDvmAL/x4zUA2wVDToXdEyWorQs9A8Tr6jcNNLCive2TDuO/q3F4IhYNkGat9adZwg0rD4sh0a
6tMH/UZ/K750alPiAsZZZMMhDdzbrvP/RMEx2/zyhyTatULqeUzYZOweI9omX9dbfRHqxG11UJEe
rOJQPp4PvlyxxKwjnvsZ87CN4py8647LxX7By+/ooa0gSYNfHZnuLbNjJt0m78UZcTKl7cdBy2xk
Rg2Rv1jzoc039YGPkz+pMEwtdrxrmVEojQ5Yh+MsnIafAjnQtP2Re6SIoHAk4ohCMxjfSeXd6ops
7S6H4nFdcxn2DpXeWngNXjHBDK6goNKHo3M1rFW7OqjWprZ58QtwLDNYJkyoTHtJwkMIlTin+IH6
ZZNtsPT5u2V5mxg5zWzrVKgtgMUY3esSVttH4eqlU0NQKeFw2+fI7HYFthlbGKsKOVGfJJbC/ahA
gu1rxdJsNOXZwBLDzIY6eLML09TYPlaqJddng6Ge64OI9PCtimD0ndZyqe9PeDHIWlguGK2yOErd
9b1er49zu0R0aYu5KvGcCT7Yic5p2TfjDBgWN5jh0hcxkXMwWlAjfpkDv/e+dFWblsuX9kPWJZq2
FFGtTkAHufJgdw8jC8Sug1d9dCqzqxj5IMg7dt/rwwHnjVn3d8xTcPqyDvjtkzLBHd9unBlZr/lO
hO9RUR2y8og/88Khfy02YnFE/0v17+L0yBpAmUr1PI5l11nwN1VIk8ycNTEl+SrMqz3aLd8HS9Pi
rjuwswiHv6cix868uu10tOnNBk+9zu8C4pcjsrfNbA4SBvVdRtqTDkdE6iRTOY9nOD7uKJtUgdDj
Ovn9pvVbUcfIuDIlaBvUYqFQ0bf+u1uCOB1WEuQ/am6omILeg54gcibGgOXSXDfbKb+fEmtpsVIg
FYj6DN29XAM9CDTf3LwA2BHv5QzME8ogloSUkNI81rI4SfNzFLWk07fTJGNy3/a+r5EUZTWEWXIz
skbsydZZJhiKG2kgCuXz6zs2JSXUe7KOvWEHIusHMj+Ou2WQ/n8ivCKtJuKhZtEl1ENRGeSfiA7u
4AGaVBRz3/bSc6VZxeUHaW0h6ayE3Uf8g0FYq+5aSHTK1i482Oe8cccETJ+Ohw4e+XSai85if4sr
QaaMZwwjU6dJwbSeS3dCTNJWRLfcMGaSS5YknSpjBAP63X3EHmgfCw4EjJTBga2Oa3HmdXvZvHWR
uzA5dK10dsU9aQVUYbw6g4cUK3QqB+VtAuYv4c+yKmzBhDASyolI4qxdzns7ehqmblMFhUNRXvzl
jaJi0BkVU7ZvEeMJKYpZ/aAvdRh3TV9lcLD0CWJrsuIfuWjhAlN+W/L7PQRUcMjvHjdDZgHbDdNL
xC7xlH3YP9GrF3dlbRo3qL32biAYlrxiqn1Oh1wGviWi6Wpzk9SRnfHh081utSP/A+nWm9oy0Jpd
FJR6XzIlFxJxwM4Hap7H29GBUjfGvey/0F40YiIBStswrpcWoxhySBGBeqvYn8PIuVKl0oNPQRkZ
W6rH6mi9Uo9yyMZMhgqAKCuSzYhzkdHaJwJBImg8Fa6MOkKtBnwCwg/mPKQeLBK663URZni7LaX8
DpZ3/tMUSSEGuF4unyi4dHiepg+YXpa+2j3y1DkHV3Ga/U50wN2h4NswBvbpgd5Ys49Na+/zrJkg
ZERPWW7cWv/B64Ei57wvmFK/0J2Y2QyWes5p4tKHB/1HyYkaaYnQ3FxxAk6cNlvipeVHOkKBH9wg
HH5e4Q8w7VTAFLYUVhZonK9hftm2B63bPW453CS3S0OamDakCPNGmG0E//o/s74c++O/XNzSUaqY
3IK4HBXlKwKV//YddQXWluItW0z8+W6MXXGT/Kl2vpvvoKRvwMfcb2qSmBl0oOmDiq5i3jhfIKBM
QNMncCB0QMiejBGcC6COKTqZ/3UU8R7M72wNBQLJyRNdDMxAGCXXKTx3gRmSJaS+eflBPvmNZWhC
oK7ZG2SPvwd6JgiMTsjjkXPImFjn6EAXEnsth1ro9oDpdrsbQWlH6qDdD99CvJx2DrTj7dw1oZhy
wl5B6OW+2mdRrOJ+yP9PD/fn+4YFXxkqStGo/dfKWmbAD5vubnbhVLRw5treSD+HVTQMt3Ux8BUR
wfloqI3DIMm2MEhrP4+v/GuhqRJ4KJZPeWd/77FEuaJ8pefRdAoBN0P6IPU1gmJmklbo2Wm7fdvE
KcOpxnLyoutElRz0DnnXj5XDIHiMqP2J/sC9iLBCxAgMcopRx30xO+ihsgsB9c5yAjnLa3BSLIrQ
AZHwJB/DnhEBvNXewuBsk9xO0I8qjZ5YsjIAmVqvYWq5cYAQK96QM44jOcWkjAtElRp0erQM+RU3
DUZZXsSu0u4Rov4t4CWD+Np4tmVmKy7EIXG2TE992REFfodmZDmDVV/QqbSJ4ZhQRDjmhzl9pjae
0hydb1p8VH2lKaPMZheuDiyUNedjU/INZG2/lyl1n8U1lYU9onjx6NiTk+i61GoVXkStQrRXX3Zr
uPLWLfrRRGwKZHnyLBL3dbbT9J5ll1qurBBVGkkdmRRQlpmVSjmYbxWW1hKtWB7TlIxmkhLVPof8
nCK1S23/QUQ642dKwOxiLkbi1x8phI8Vn+/vO5YbuoU2pr4PmwXqZpEDR2DXNGJknSaonQoTkoR5
BImnk+D7KP/QrnkvcdWsfdIoq5EYPnISxKVA73ARGC2aeAj0ayLW08ZLGR0oN2yDcge2ZFqSK/ue
QpxvXiwwbpN8p/a7hqedYoI3WhlgxOUCc3kDP2DRIkVEusm3dxpteMrqPkHbAQAA/P8Jq/TZV3iM
BucSFZ2of9UJBPpgCmHdXpN4XE15xVUYBnv2NkqDp9KPGFUV8kgh4LFaRriqXcajWRps1KM80t/s
eHpYoa80svURY85T1p1zPCmIKRe4xa7ykLdNcFSQykefGwEJ/8EWBzO9U90dxDAb3Yl5RF/f5rzu
Mwhlx0S2/gAPP1TAMNwkEQ1ubfkXYDwFV4lbgvClXIsjdIs2Ep6GAmdpHevf6Llgh23zCiIjoOuA
qUAT7cIDZ1Eas5aqri41Qm08TDwrdLl4OHRvfG2qaBYZENCBjX3AksF7IVO8EJotoaOk/E6OnrKM
ke+mDq9VPwZ9Jb5eSFKxDHe8EidvQ9GEEcjrBTlBHD8Z4QS9n86Hf2UD4R3LSP2TPIkyi5WlKWdY
0knYnINYm0+9Utut/ATYDJN6amLyjuFsQ8KDygLTP3yrd+loJtruOmbOP/qZzVLw5Se1PdWEovz6
IystZw0WeOrrDJTGnn5DSYeLYJhZLOLHLKSD6dM+RX6WQ8Zlnt7D65S7Gi6ubjghUSALqHkeN4Xb
a3ebWknjOD81+ezOqpDTQiUapN8HRsqFZzIVvlLwMP5LuWVOYProPO4wM64h0BygRKLRaMz5u/u2
kVb17/2eb52wbgjJUlYOFv82QxXKbEGv1dbm6Ws6Luwg9UYf5J6DDrHfpM+9+9ptlnzLFp9Tyfsy
QViiP65uxjX8Qdu6aZQZfG2gfTHkxdykzEslc/6YmuDQR2TpAdBrn3SBXmQ94uHj94+4TR2vOFjV
PJen0RXP/MeaLe89qpRcsWxtq5YwNZESDrd83eGeb/Of1U0l4jmWMSUQxrr8dAGHP14cH+4Eg5FC
tVp0n8OGUY6MBAKVDKO+NRvXQZQsAfpqCP3I5IX+3QyH9vieIfgbOFkYl4Rm/6C8oCKhhoFk0V3Q
KGhj1jhUmk8kB8NEJcBOi6DNjQOPVvcF5LvuPGj3SOgyIOsPHyQ5LO9ohwefCCwi+ksWoRhTE5cf
92I+niFGNCUoCtIldztfNDR8Q6tYJvmGUwtGi0ao2mEUxXQ4n2qymAboZza6+tSPNUAaTtDOtTB9
koRHJEVR14L6fTn2PrHZURsa44Wwp3iySa9NWwY8KDBa/YvdG2Yt1ZhL8a7RRSLNIe4oTEedeD6e
s/tbsH28WFQ1CT637XLH2W7RaUxX4nxeHpbL1FWbVCrOnLPjLa91YUed9dLTkZfjdzKazZ7GKpue
MkPzRZgForOx76pf2NsC/9pkeQjUo41fc67LHz/2avYsX1OtDRyCzRf/FxmFrgFtpMXuTxqljsqE
yno0gJzeOYOWJsDXlpctutdPytaAlAxg6YKtK0+/R2vl8XWe1AWElk6PgNrDjr1nbKbu09SExXM3
peMn73zmhgGUHYp+Ko/qB6VxPN8LAzodmD1Ct1SSgx07WFZhKN7+/HZZ+F4g/uq7mBK/KXJvTVa1
AgXC5c1ii9e73FF5DcToksXcE7NnicxzfCuVECzf5c5dpmYIwaniMREnoh7H6zubeuMTGclnbrdO
xA242Ad3Pm1rS23+apuw+u6n+pz6hbwnDE94DAvXkgSu78WE/rCiJ+wv9Wbp/0udl3yZEjr+X1zQ
wM0E4pmu8W1eGIx3PmgK/SGxrtN5bJTOFHTwTJJD3DM4C0XAfQe3oOmhc7hvy23+FGUEpLM+lgKA
0JB9WOe83xPQYl4nl2P8kuGm9DjfqQyZ4o6e0TxGBDINjroK6YZf9tB8d/xYpb+zVcYvJS5UlTWo
VL3LAyZTNiESEp+fZZSjp+21+Sj8N5okRd1+FflZxpqOyITb6wHPOezoWlB1wCDVqMkqptuhuz/c
1/YVpBvE27yP9bPDc3+sfdUoWagVF9Z5g7Vg5Ry547xyFgSCRBNFyA7d/sTZ6GlH9yay7Yuev8NQ
1JJM+B+WAE/TsLAD/K+8BHYWz/OZnnrRsRrNZWEPIPSshSTnbT3xJWr5jOknIvgsp/uX3bSAvu1n
3oOPlF4yLxPI8OwAFYWWLjRJ14BCmlh6EK360b+OSpfWLTb5WqZCQdeAoSdKKNepAx41gQWHK2X2
eqIZvxYnFPEwJ/HT03y5OyaYQ0gC98N5RzVUsa5Il8lj+VTmzWN+5EIEOKBYYgq8Isg3cafXj4M8
y629kQh0sqqcX47I2uJXnGZgPsFBauHbQhO0HMD5LXe9dTi3OVDVu7f5Lb6la/ENb2ShYoGL1LNq
bdSxejsO/MLsP4n3xd8d/4ejHr1MGOAOzxG+xGFWFVDbv9rD8mR1yVExtnWcilnyZxo9nVix0dQF
zUk5DtHWy48yio2x7971zIiiPqoMexFMeEXSrHjz58H5qF8ZYRcTNtT1BYjttZMfhRUN+lYymOo8
a8xCLp5BR6gKwr+EoIKFM/UiLoUsRo+dghtlz5h9jvTqm/4RmZg6wX/2lU7onwWOn3/gxp15aXSV
kNgn++jm33wis1nZNic1Mc2GBc4sVhpajvDnkoZ+qaxGMSravM78N6bWPziHz2GAXH0qbyD9H7Ks
rEo30YxlQ/vAzZj7Eg95IOEeuH76qJR2cOAwxigpfvdrN+A/Mx9qAJzbY2uzRh8z+dNgsEoVLx0y
KnDh16n0y/h+KMN7PRVU2/DAM7qgXslqZGJTnO8Lokp+BMj2SNud0NewZ040u2xHL8BANL8mNrn0
i0zncEr1cuIjqB1ez9AAIJhfCVsAfxloDHc3aH6wPaiL57g4UX0tTNdv6Rbzry1qbEn8ZYBQ3iz9
0or9WKrLKRhEG0s1X3eu4zPbYUZvjnOmIfnkdptceJPDa13LGghvEJtjoH+v1JYIYhVp4wfKywtj
rOz3O5qqGyPjr6UN4L1FBS6OIHQXZ3ByA/pfXmNqbNlsmpi1E5hn95oBYCRbw8cUZbuorfLUdei8
E9CQuJDMnxS4LDhtRGt5Uo0JTKLWbvmPNvA9C1mAHtydz5dp8skdYlw58FIqhZtA+oySFL+NzOH/
Yo2BiMtfgtUDsQO/N2Ny/TCkQC5QVR6eTw1Xn994YKSW1EbIWPizxEZN4k4USPpwH0+SWtklXg/E
wJkrZRkTwLgOTWsGVz1Xv/zxU2V9dQ3ZRF4PbJZm3DZ1tnGlmUud2h/sJW92GBXEltcjJrYyN+jw
EFq+Tl8dzQrvDTJkAw7BOJ3G/+579YjCkSWzUSXSbbHc35B4O42Cica7Qr1GYV71BBAaOHhdwCz8
L6A6nVMydA3MvXX6/HP5/WrsZAT9EB7KK4BX3k3Oi8UvVwOA8FQRz2l9WG5fo/uzF56ajAjmWTE8
U2kVRvlaX5I91gRFIc3Db82ZwJUWkLwf+WZDd8oa6LZdh39/l/AZYhfoGe/6OIavtXbH18jv5+5+
cylfxV06fnfF0xxx8XvrdhvqWG+hEPSdF+1RW8no03oOkdWryId+RB8m2MsEn1Lja0rnvYDC/F2x
Bq85arI+oJ9C7LWahX1MNOku0yFfiPuZZJky0lRV6HZU+Izgl8dAuSbgaGlNtr1tbhPgGqXwafFw
eYV0QFBqg3BAXvJzCsWR7wmMKJGErIAKvOE+ZleqRGRx1slc98r7PFPNbmRNgn3cDymHYWuJiqJg
cq5JBxZq3sJpVRvKpJF5oDGJSaQ/ISQ2mLxA01oMq6csGBxiWnXA6YEJNT9TBH/oZYIIMAmfjg2B
EyoiVARnfI8pFogB96du1isO/Wo7OLRPwuwCl11jh3BVtu3XCzW0gsbjaMHoZ7u1JVsQ8zeBwDtY
Xgn4F+1QvWVn3ksi4pafGuTAakVm6wCVyTnqkahu2Q9eZiNyRKiCuWtvjRNoO9rzjGeFuoWPqeqh
nxEfa3EDpwiHE0Lb1BhLStbldNy9y+HOzeXYrrNJE7R20flcgRxZ7VFk+voDsLCMXonvBbGXr3nz
NltDmXAgs8BV+N04K0tpxrkA14K1aBi1uWq2LBX23Boa4Uh8qNyM1ksF2Kd9NfWPP6LW232jh3HU
dgedkc5k4v2BI7d0WT6b4/tzFWyIMOUdYKJeLFuvoCqiqRQQA+3lxpNqiSW4pzGf/wlLaogcNMms
E8RKaSPYyWJpIkP9G2fGbQXseaeCYAwXEFIScltGkgjhOv2FFvjs3PxVm9yaxeH/6bUzuQmZtVZL
iTAigyVZULIieXPb+9zuprd/PN2L/x2qubwWxvQP/Do0t/fYz9r0QguIVCwDhbF3VzOTJo7Aalnd
nZt/APAruJ9J5s/4Hn8SPe2dLkVKuQnmvVQ4dpYEETbb47Ap1WVlw9OyKpDCSuToVYys54oB4CvT
ClCm2yTpEXnwV7/jo8bEgUQvyt5hLolOZMhT+UU/3OYyJElLkCUpIesMkRWdEaICaOSdfd98Yp54
4oRg2xWdyDbIZfDQ2ngSvB/YpORYOGziWdKojRXAbHWJe6nhNETc+XUjhnkwpj0mJ7gqBdMeazU/
hqGGnnvm7VSLuPGUgPju7m87X1Hnl8Olj3v/2+NBtRSdnsQN9WCq6wB+31hgmMXtLQVsFv2W+3CK
ThuoRTiObiM3ZLbUv/VNkUCDYDDD7uwlVeMZxvVscV8fjcJw8z3sSL6OLBFWbtnww0yz2KU+jHvs
glr+6L1Zdkkyvie5Yk6I3M4hM5ejQIT0+0wtVRppxqdEGdf7nrBkZRcSC77WgfOa/8eJErZuekfN
dbnv8/VFbeZ4fUJ4pqw++Ou9ppAapN7noRGAVBeYSIPjYm/1s7ddrPMTdp4d5VbxT2KaaRnjuTzT
Zr8kAK7s1tQkH4SGlbfEHIE/DdhH1C7z0/AD7N5ZlbsOw2wBKwMkvwFW8Py4VtOIT5Fvar2vFcbX
xf/Q04IEhxSfBJ0KB4i2dDvyMzIXIYE6AKJNrXY8X51X/eQAzW3pVv+Xc1+obIDWC+QMl6FDT/h9
g/lkGJhH6ma95+aZakiO5YF/joD+1pE8F9BIABtSgGQDoFEbr3Nb5OAevBLTDaBlop43V025ho08
G/BChiMOz/R2vLOTjxh8ZwPVsvdrpi10AWcrXTP/JmTAJNqgygMei1N92LyBVGbZfa7zKqxJyCRO
xy0YZHf7+B6frkZnZhZaYIynMju+MD8LAz/kpDhWHmlE2F5DWaFYo2sMoHrwXCX9CoEnjUob6Avq
vv6CmiarXreTaNnYVDbIZLiINTtO+VHqQrDG8pXjBzxSjmth6BDLZVBWhv0oP9s5g/XD2dlfHPuu
ELaOMuh+BpfNe89VzWgDZu9bF9cGLrMbtbLNerhxTOlt8Dh3+aIaosqRJxRe4FMLPXJhQtx/+L6p
dgsO210xGx/8+pcOUjeIkBnT241uZmpBi9spH3blfHUlGTQJDcay5Yfw4gWUAhH7kS4T8eMRVFSU
uV2x/eZQhqd+aQ2sXinBW/sIuc1Rm/+efePvc3K0a+J219BUhLidUI3gU2jDsHvTMoxhpj7VL8eO
9ZvWpFZrGTyjE76IrWbwcR9Nlf83AeT8qMVlQUY3H2I5+0MdBGmx+/CeC8M692AqIrkUoBwcRLtj
iU9g/zqw5pG7L6NtnqeEeNmLuU8G/LwQRU/ighgmEd6K7X2g6As4eeQve+uXedoeOcuteRUjBl4U
9usbD9iQo6Yy/VOrwOPmfWDu4djUhFL8Y5MSnnDWaKarPubJJWzbUbEl4k2528pybocqy8VCaFSF
AxKC+dRzZUJVrPY6Ox1NfJtd69UfWZOV+K0JqzdMF2CUmnbolS4sT8zOhwqwnUAFE+2z7p+ZK8tz
IE13uJgrPr5ZGeBhcyLGR2lkUOjIydlDkzanmcblRiKOT3Tj1WEGds0z2EL81p4X7c4z8+xU5atm
0ajQUnAJf6naYe7mGNZwul160xnWsW4/kXVPR1JCLYZBtvQ6V2T4clw2SfVtt1uKYnnls+eMLcUR
SOyqD8Kkf4nms3oozXAasxCoGPjYrAGDtVgWAE5p8+lyvaDG4IuAlp7GusZwQEPp+xM34tP68pOS
Aor+SnmJDiJbm/PpceUmJWalvne1KPTRe5JVsdB9M6Q5nrjV4A2nB3uPTOa44uvz8VOYHXC59EYd
bekuzZoVpKc2LSl8hdlx8koo3LYP7MP/LUU7g+1Kv+NmYNYsrVlXt3zh06r3W8yGmQ3uyNfE1C1Y
noVfQ0z6wdUKJcJsutyueTwaesRd0RUc0g3bKUZyd/iuDXmKkRGS9SsaKeQpuVrvcodqSzqN08Qs
AodOWpL7jy8o80qkD37Ts/OsfPbp771qQXQKsBzBu+StJaxke6TDjJb4Hk6Jg7mZbuQiHCaLGTdw
Sw1zbsfMXAEYRlxgGk3hgZR4XO80SiP76SYux6Z6JGvMunRaUfnHLlIe9lxKtEmLJlKY4vmlKkqy
zkOZKPIZxzUGE4x/BTphO3FVmpOebNTcgUWIZKt8wkZf/7Qsp+Ao4syMbOP6l1s075WwwZe9wFWG
6/ztC1bTBYc6CWFcygcB4RhElM6RlNg9dmrTbR1h7bFyO66FzINFROXI4ejQT+WHwsMkpYzIp2hR
LSZjmI+eaH/km4FBNqI5RtJdsZiICF6GrzODHnAI4ANDP0mVOWbi/c+JSSLBQj5U9VwOUhSw7S/H
NklXivJI2LMOEg4nOML/FD9GQHfdyJlQpzaBmaGU9qCYKYAUlJ1yDtaW/T14kT7n1qbwMR07i9D/
UbTpfbeBUG2CeZOX/F1Wn4o8J3ZKNhyZmA3nvKz5fMVzgOSj9wveGOPhaqITIt39dPrNTpsB4qsO
SyoHUZIV4tFmIMC8ZIGGo8kCjuNeVfEqPYHKRaMZmPFsfoct8FwuLAYn2Z58VRp9ebNgXifZbM+C
/8/vrNiTp1NoXGRqNkf+nz72TrCsRYKI7EntCaFUX8pIw0TNS8grC1/3qIhWzmQsUrWlVpxHS9+a
vYiUPuW5YLRdLFx8lb+N6GaWrhM2b0AfIdXrnfigaRu+Q/5dh4FoEPWrFGQXAHlRJ4ANvZm+oUNA
RhdZwJZ4dFCdKC12kFMLOY225GBFstTGNwT/GNQL5iNnzJOmVqIXuYnWxtqReF/H1yTApLJRgbc8
rQk1Dp0BWhV2AeprhM3mfXQDPOajMO1I3ncI2T351YTvadRfICfVPg2nlONAEUzMuwTDtl8pO2Hh
J9Khow1/W8d8Av2HdU6Dc91B5GJazFpD5qI9n4/gl7pb3NaRvYMbukgrHrpfspInMHbingDAWHGv
lKbNmkXflisWstkFYTuJjXAnYnELgaVUeM7jyolQOp06okVZk8b9XhFjD1OCmBIXuVGkecWPD0KJ
GDujEFLyamNZOJHuLrMPVT89vXJJs9cxDuYum4xROxaOJvh8Z1FoLdmZ3YjS53dKgoPZ4aaNAmxO
e0qHvxUt++sfQD1HAc1wIgx8wj3B71hWoEJCQYXZgZQpgcUNn/cX4cK/L/fk1oFpQjfGmvD9FBzn
V/Bf+ZNNWNS80aoWndQeKJcist1Zhp4IqU4e6ukwZaoSDfgHitn3dpC2N12h1vmcWDQffYwx+hsw
sa5DSkttJjM7dth2MD8AZJJyAtV/oUUydV7JYEfz0f4WDwGlNjN1trsGN7IGtL7d8GhNt64w+PDe
XuKYwZ9QkJFFrC8bsLP7I4RK9OjU2+xlV0PsA9daeXeAqoIjKptrCYyLp8xAj/ujiN8yvSRp8khP
V1Ju8yy/6ci3bHdn9RJ2LbGqijOy2tfBcb7C3+2zL/Bg90uO+GKfA2gDVl6ebRq3joEveWeU9lJ7
RA+Q7kasQ89U/y6g/zJqWbWwB/+MBkFxaPuXr11XMaL3OWHT6wEm5U/o9UAj6COT1fNiZf/puhFG
yzQ1iauyqU05pdmJyGplOCNGsR6kZW1bL6uG0nfHcWY3x/gzg8OZE6wSpAUTF1Z3EOVnvn96JQIy
++KdedMxt0IrUev5gbsGvAR8ymyumJ5PyUMpXX/rfhINhsxFyjeiRsjHBbyzUsHezcPN3MOn31NR
s/D6UQcFANBzUEvEf+0ovPHdvEkvJVpi4cM92MuqrEfL/+qtbV3k0/TNwf2vudBpIJkTckQmVXpk
b2Q/DNFWyRqL9uuZ6LY4PEBoL9zbRVQtlay9Qb+F6RC6t5Rrq67zK4CVcGGkZDPR8zTKATNdLoEU
Gnbvj9qLPlB5IQgYiZpbwDHjyCjbnkI8moPn4+9ZO3k/DG5uGTAwgSuAwetuW7lXSf9wVEx65MIt
QWyg1X8Z2oKCIVV9RhGX2uEQ4gBau+F/IHV0Y/o73qS9520nhg7yxOZBIfUsy2K5B2LnLum/Wn5V
aNABcjow5I9/vFKYU/ks4H1H48v4D35tp9SRES9zPJaCK8FNU8F0YSY9ffYqsGaKTKPGG2oX4Zn4
x1BDm1qruLbB6jlBGJDOe+PcnBdOpiSP3aOnXtjF+pI+BXOnBTjJHFI0g220XiW9w5oA2gSXUgWj
CQFhDQQ3WXTW/ltCJgFdSbRqIXzIgVyjc+BqdsOCUiRn78L6qye/JYu+beeDD7+yEKtltuyEZb/g
bb64oV8YGUfgoH5AKm9jNZWOzdBNB40iYWrw9nD+7VYgoEiRu5c6L+VTvX0Qk8axq3k8NJN1LkAm
CvT0WONImkcuy0lMZaZ+bHw1PmSRjyOs1ATBVWXYxrkdbAN9haO83lWrjKTmcb5CuOhP4tYcUrdy
CiqM0hZmK2ZUaR0Jf5VuOMFBFkKRGJ3/hULNmEvCaiVAauA8agXb108Bs1eCM6rlfnH0dppUMTcu
+fBve1+cxISfOR0XLnjkVbVvMoBeRU/0EYFYnuEUg8btEexU4HZXACdE/jdtMWtPj9ugwvrYWVaj
M2QsfXEkkPMIwdZjzDuc/WnbHNMvXxMUp8BAmq+XsVPUda4jLdcrTTHkcK8Rjt3GU9kUTE+p6qCT
ORLYdKSps2hrSO4RA0TQQh/zNEqTvwMa3g4JQGRosnk3c2MSaKHTPAcAoXEcfSaiyMub5XM6gk+b
Av1aULTVgBEevUfFdM+OQd/J4nHFRRDRmyunLvPoS9Ar95mUhSk13GRYayZHm9vnz1i3kH2kQ4qp
/YLjpvLh7KMx+gPfQGwNb5ta6+NZpq4CSfYi7nfjNTyAThFX4SJaAQ0xpopWqkjahaw32DG4l0E/
2HnSx7FF98C6peI5hJ/4KWM5XNJC0hq58oObvZQmb9Bc7CW54Ci7aK33IDNEgUUu8lO4QZxVK9AX
upHjc8qIEG+0vdaHtq8iKsYSyfF1y5z0SOucRiagbzesOmYyRo03A3viP9xRW6eWozUIR6ZmwvQP
KcIuSuXtiCTLFJI6lfPo61hcnnYb4+DN98VzTYnOG6PcvDEXbrIoFWBmSDWVpWclSu4zpn7cnGXp
kB3hFrYsvZkpTYMn/5A5DuuylqBrlmwD3fuRstEXT0PwPzggzvkJ+wlsRq/jSBYE35Gu4iPgJMS1
3jDVW+SfwwzIMA0cThyXyP0GMcMeMXwIGApaDjVwjEX3XyKx0nd8SdOGwOwvoEcy8KPZbcx2pMSB
luoQiaOC4ssfVpDtKPW86ciQSBVuOt9H7sK9S9irAAAitKDLzwaVAQK6i42x8m7V6PbuFolsFZ2Y
/QA2AzWgJgrLKPHIhvCyrE6Pc3lER5uSZdGu4HSjbZXMU7mhKE6RgJQlVePrWvon3h2RyPDpOt71
3PDbagtqMq2BO77kjZGaG/7phcSJ6isnpuo7MNrNYUcU20Hd1GT3NQZ5t1Yw1T1xQYBknq6gQvel
GBL4cyC5DF/uIxd7tP80jetfx7uQNEAua6uiqAWcxY6MMWME8pdQ9wlmbc78MK9oRkBc1Qgn9ihE
5RC36c/MRynWarziq3lfNu5EVNRfsOvS4hDxa+F6VBEr+Flh4zO7x1dJ1K7eSxz65PIwchPVpdxh
EKneT7ms3E1nRoFOe2mwvRYLiG9PRWt4FhKCw4yY3HSXxJnMPqSg1EnUlvVchkqHjGrQ1u94P8Op
Um5t/zCSikB0eHezCkdnMb2GWFxq8S+ZRkoOPrkFlLIDpjm+kGHW54OfEWw2zjiXxkGf2AMdfjE6
+LDwmRpGogxC81kwLHu1eYOCCl4nV0vNRY46R1f/28PzqCDO5yj956Q8Va38Pa4vIfaT3P6QqAto
+WzBXA+pSmXqd34bPIlbsgGRlb1hXmIzg3q8HHQWIgTC3vPtSd7IDuOdWBLYrxLSh9EwZnhMTH9n
UC0d2XbZm84PLkeaPgcz9cQF07kVoCCM+DY5yKUHvvtz8FoyETBxZotzU2lSWFBMkOa0zIKhhdri
TY/5VX4o54HEuDR78Mu7g0o9/GFsCeKvBQvsYa/9usRSaFb5T/Sr5OHNVROvjUFz2ALkXEPwgb+0
+hyFlvBDPQQYyliiyiOv9v9s7Dy7yZnwfH/eGIp1rHrowutpawJd2uYUp0bhRsNZ6fKlslNti8+F
d9cMlbqINs5K0eRf+PFWJ2EwQo3wmm1ZMEVUm3+CyrQuHexqVq/BtUlsyfdpD5vObtu81et5ir+i
l0aPKIl9Cs3OX5HvVbPNCQanVvi6YYhx7bMn0Q6moJb1pOn5/y7yZd3TwN4mYFThfFgi+1ocSiAc
NO8ZC/lWnI3w/FAm0zyUDvB6oK5zu6+pf0mWG4WXCFgg7UCeWc2vsH8Zq/ipO9fJcRC8A8NAMU/i
5kxdTIocXMwhz/U8qsr1nlUHqiCRNbXG0aAHa0fnG92QrhxTmbC/l/3WxOkngEW+TP9mPlKqM+99
Svfa4W1SneCi7xw6A7x60yT6oL+gIUoX2uQg/U/H+idGX4yphCRI22yGt0AwQiAGQkir5q4IaNTd
VZXN8gkD0fSDsxIGC9wxlORaP9LeCfuYfOmlSlaj1ZpOVxWEsDF+ubeXjMIj8nwkiTjpctScDxz0
8F47EwPsW8v/SrdBSxjHIo2TPVLs4AnI2QtFjLefb1jlCkC1Ok8AULoazjqzaZZ/juAysK11FxZQ
gEGwK95mITDJiQph3hIKhb6npDeZuqDjJ4hLHNp/Q/t7e+4hHmkMewYw/Dr/BxagifM3Y8ZNqqow
K7l8qV0SpQcOrUUHVZ9QOGtZZUjOL1EueJP2P9htsgxQq3OLS9q75ArX2GKPspH5WVAZC/Uctx7q
XVR8IqKP9UUkj5Rz/fiIuHL4pOEt5wbjnVa+CAcNP6nMoZiQ6HV99ZyrOI5c0ma/36zM4fiOoT8t
VTyXfrjcUtxJnq6mJNi1RuxRsfbK9UNWpc8rSpH2z7FXC0VJKEjlMl56lcFcolrd3ndvFvBCnjOU
tNz8SAruRC3DZ8JX2mVHfgbedMo1wa63w3vcENmpTEOj2owAiz2IcuZL9qHO8RrWuxNjk5tHD0Og
eOc98s5uy6P85Rz0vfnbrxAlXhxXL2F5ApiQFLeUZ/CbHQe5+dlpitHuq+pDuEDjneUhXQE8LdaR
CL/fr+6LwNs6pbQLHaNCzndaY47/U8CJOPRG5TDuIiWWPNzuSPi3Ui4QrbE6LoynT4cIkWgn/4s2
Gl9yjDjaQGTRFLAeKRpUTCDIB12ZRTwH8VqnTboYbzHAxllzydUtW80VMIDQwmdJy4iNcboycXLd
V9+EnFnhvvqPeQLzIZruuIoMR5kgXenBnkrpz4386doQtrhdt64ZOwDBmUNUGRiQi13yvtxDLd+K
fqaBhlsgm3RDwqCsvuSUy5c3Rq8FwqhoBDHcSOpey9ytHUShkbX9uHFqhlNa5k3wKq6vHFl42SaI
UXRh+1DUP/s2SNmZTBcaqvHm8LZeEFL165uIHZAcNwioa4h8KYrDDXqStZQuET6X//rCI/eZY3P2
OVVFlfG3kqDa1HVQbMiqaRYW/i0t30ElaszWW5Zx7HdQWgZQjXQ25ETQfWg0pBdTJjFvcRPgGXU8
NVbhTgQCezHQKyaoxm7Umc7XDwQFgE5hKXoxBSjzpI6eM2f1aoc9uClIGBo6jqzcfv40yYJ6G9qb
9UllEurYRfqMemjO/81HZM8EuQ3wxYCmTOMZ/v+gLUG21YKDWoba/tuD5W7gUWYvu87xj7ynCQ70
HZ/lTAgwHICGAdt90zMnwWcbjdvTU/m5Yk17aAtVX//DedaCwUHp0/VPsyFZhFQfmDcC+kOwQ5iO
8PNVWFK8pxEf7IpF3RMWo68mNctXWJo5bUhLTkg0Pbw+KrK47xPIm5z5RiH5kcrHDmiaccO6p9MM
i+epdV+RksBPlAaf2ow3moV9NwGgWQRo/ZGtiNPOB/8Ud6G4KCUrbQAOwXsUb4zBa3ad+T2TO13U
r52T8DusjeZrNeXs7PYaUter9EPSEnVy8Kc6AoNoOcTZ4DGNSE2rh6BlSAKM27wNeZ1hbxN8rZJb
9VoT2KmNyVduURO/X4SB63IO9wB5WGUC7tN99n5aS4VvhlTnu8GVTLcG/hirwwo6FWnqFxUOu7m2
s/ykt3mq55Xv3RJk23FXqsYcfO5R4IcDeNERu9ATyNjPK7luuothZis2v01iGswDTKF5EXBJPklr
EO4PKRhiNTLNd1nmwYb7onbZujWPcknlyyi/kD6b+bOibHpQpdq/vGeY75B7cBfXrZ95Aq3xVXbv
Q6xuR36zyAfW72G4mCB0S16uN0vdmoFyFoQ/ztVDsTeFh7NQwcw5/LXasztVXOiIuMhElEuv8NJ2
aiCTBzv6aOF0RT8YbjW/ImA40zdH4DjyAQIKAqyw70CzJmdfioKP4TPas5D0fTKNKlq80BxxbNSB
esn4fgq2khvhxR4TRhuJjW2B18B4dwgqYlhmyXZSN/0/sUnSxOweB/TUpo90cw6KAkydE+M3RLWT
C3VcfagdwOb5BtpqJdfcxVjepFMEGAGO3gqY8AAIQ82Qyu5msKrwrsWDqy1Z2T5NYkZuiqL/5kCP
4OS9pD0ApdKLOsP9PAA6IPt8R16etSX7EM+gcL+FWxSU8SgSX7ts/CpBcR2uqnuRHmpWLTFMEVx0
AO1z4jXCMsohsDof4KK5eLdCJ0m3binK9UkfjYkLXLzfB3TK7ocJO6gRViOdcatIuGVDQz3W2ctP
lLTOpIkrxlKxVP2TXzjKjwldcdJUMO2nAs6dEAKaX45gPeiNLO/ZF31LoddpCW3Ml3MYf8QIwVYE
CcfUUeUl3z+unkNE+LoLjoKL8U7J/R7UoujmiGnuZWRtTmU3YvRhjB1Oiuv4648G5qflr3X/Kl/m
G3yXVINuOXQSOkLDdtIKKbiAk1F09n/aGau/cdG8h0pV6cHQlW/kBu0VHTiZxzoLJR/BTn22JqAL
kfb8bAjJSeYoWvZQzg7auZpo27o263ONC94/JZttEbLdu6xTX00nSpi69REqrb+BEmzHTqZX+qix
hUWdXtxsj1oGmIIQTlD6F1BpGtKTgc2SYoSvPcyF1XcrAs9qvddW3+xdtvAc7/jvd6H0MP2Jq+qe
Rz9X6wrPiVnMhs/NGO24RbDVle42J20O1Dhdv7tUoNy5vAHPKjhmnwiycsIQRnDlD1dK9wK+rR51
oqE1Td8wORuXXUA2CatC8pEcDjhmFh98atLFUEJaAJbFYswtJJksWg5Hh6rFmzDsGNzv1nR9n5p6
dujiu1WXI6ehpdgwBZxkD8k+SlGJifi25rt4fSnqfB8sOf3xnJ/xNKiEWvomQUVGz7xObkllT0iO
lo3KitGRYFSVIxlFYtgJqR/frq5vVorJj8upC3HIcft+iXdEZShTSyyRhHpcW5T6ksddJY97BTW1
gDGP7C4RPxi02Y3/bXxl3tfvQc+2hLxiWisIgqLWh0ITbK2lNmOg8Ld2aISpH28slnIugQNNE9WW
QBodRbUZ1ToSnpwAmz4BR7kyslD9IEXT0NlOxNvVSK4GeNuMa/Ni33QAqHUtVIjpS/vK/QanP2Uy
gjf8W1mijQvKRP8WPls1liXkXGznZ2UWe3YODsiNw2TCkCc/TnvhkgH4/wixBEBsUxj+L+6HkKb+
94We75zF/URn1zzbeKjN0u1fOaWV1EtcwlITXE/aRrcJGGK+QTt6zvjw+g0EvQx7Tg7N7biHUAr1
lJcx5z4PcegL91+dEzbVIpu+TMnMfinZ6MeJz1SZVSxksxMtLupO7VdPhXxwN2TDythpVKQ0PdjG
vDgMW9yPtuwfJg9lteR4xNeoALUWq7o/D8e8XsPujN/VEsXqoQXl+JbkDbpye+vdeF0kGYEbCTaU
FQzDFiDZcUp80eR53OeC5suJOtue4Y9EPj1jFil7g0sodYXtQho90kAXPhEl/FjHh6DiK7QEDln9
qY0lmJXrZRn4JAcv2+iaKOah9uOGo1iocwyvB0xtUv8ZAK1+TOzR/jmVdyNOavEEcFPgq/t711Iu
x6igQu/mNDYzyIlnkbiJyTkCa/jgMp2PPWrlVaXUB+efRO9UMxN9vh8dp4yiqaTQ3CP4vnwPzQtP
h5dldYPmNiAB+haQcPW08N1tsktMAVjic2xRxZEMsbkHEvZhEWWNc9KUfvIS5SkdJQ1cluCKHsMC
4930YabmRBNQSJvgfVVGigME6iMX1CIbZH4JJvftUJYY2Xqq8s3wmEt2wkcHWsTgDbSNuB44Cucp
Rb2WYhDzXV7lQU0oBcukYSPmVVKwY0KZk8bselAKRse+bwlikdqGo1HUTkR1JcnT+E1ilG/Kzyvz
0GAEhaqpikRz8rlGMwHdWg+Wku3yMvNcHCjvrXVmQ1xc+H9fRa2R/BTjKzC8QbmgiTkwhOTwhsxp
pN7mGdjHqxB0qFwftRkmkzXuPHY4OExx5LltYeEgBXgUZw2uYVXko5L4j4RJCORg9zsnNvmgZxC/
8uqfMsRI4gU5LJKY4XE7sijOrVyBHtvpQ+Vx5pANrIpSu9GZqSiyFVobkvQumrJ7dfJLcJy7FqZF
28eWNnYGOUtXZejwPaV2Wc3C88ikN7AqRtCuAf9CqCZQExuK21Q2osWLaqsE/v1QZFJju2PeQ8cD
Ie7dbMnTaS1huINPYrywDhOGIpehBZDxeHlvZkTcqqKQQOyokksI4y2TV+UPP82J1xWTRvuLNmgb
inpMhWd5bvUlOYOZLqTX1v1+WwgG1NenTcGDN/sBvyl/qwkP8Avuso7Hjy9iuJkn5gNU0y/pWe/j
1cYm7nhs1qX9DRobonxIuVa+JpZ3C6N7NyNdvJd2QPBWclW703g+B4RdE9F1jSdynQ5wKA/t1exS
nQLFmXTJCvTOEQ69ZfUvrtUkGBDyM5VJbuWeZHF5Qoq5Nx0QC7m4umYew1IuDRf4nDc/705hUh3U
fylrZYDEMv1gu/gPEl555JJCm7UMzYH7OTpJPcxBCh262WcOjICmGUdQcxQRK7b1706q0c7YhuV/
dlOyPKoKSwmDKI9JNEL76Z2CA4hCtSRuPFY7B9feKy69JsYAGXD1kagxQwQNqQvv3MR2UMxHUaUx
6J8MW+b2TA5YjoRJUooWKah8HxPZ8kySAdXaW7KZ6GhoHgteyR0vuKNxrUY2X6IIk/InonbqFNET
VsJ89EV/z1+jF6tmITSdcIx9QDVD/CqT0hMEMmsIWVopDnna3Oe5RD6b/X6Rny5892AniLg7nhXj
BD1/tRDK8Mxy4fnzZoWoRepy8am9u1Q+6q/QEU7fafQEMis50VAPYEke1O0qN9FT/ACk1xUQ4wYq
OnMt4mvwT8aubBU0SpU69+3WuP390ZnhmJpQCrNW5wfTuNR/HiUJ76umBF+neiP0zlZpcXyDDJ8k
7n63mxkr19HwfICY/tNdfwPvfY6pPU4if1LyM6ZLC3g7xY39xPhYVi6HGaN9Tx5mCsXzYO7M/l2D
ymd+kh44d0BgxkNyjUhWwepTTL0UDLU8CLd89+4TjAHbkYKLXGcI5Vkd+kEXt8xgkkXgF8BbHI5O
uas/ia9/NvUQBL9Us7uneRPfqLlQ7B+6XidAThASm8aiVyMzHnMRtt7mLM4KnaOKPJXwvaHsAZUA
qaMzo24MtpLQaQQfwr4pVKSkLg2SZPN+xtMW/5+bEuKWcUGBRs3XSlPk0t7hTBnDyGQJS+zzoCTY
H3NCbfoDk1p6SUS5vjelKIuMMb1fD/lpVovZxi0jpazZVOsFQlIYOR5hcXUYApBfKhH/Hp7BApjb
hvHZmfiO6rCz90ZHaTL5dZvsJ4BY5lI6hRdryj5dLr3cHW/o9sl3y1w8WjTUZy3TxuiCMnfccY4/
bPwrVivcdoZwJnYb8ktOGCaOMniVfJTk4cSBPAljVjCbWWs1FZlvBUtLOgE7RtztAo2pAkgpEOES
MrY2qbrTWVzPeR7RJ+uA2bgRMnQADia3WJeFml+sYJU/JsI35hhFY4y8Suz2q9Oq1fVkUw1T7d/a
oiINTYRx8ubuoC2XwtiUYozTaUWrkjwI/SM5ccUE8rGDX2HJBkwW2LT5p4GKWDTnLrQxI7AOI06H
QVRlvO0ZSakN71e5z6f4wzt9XCr7WtDaYKPc0lEpwlORDYp8XZKB3+tJVDRzzDlO/RpPYfwX8fQI
fWrx6d3zY8K97jLkwzfsqFa4AtSQDiQYbiiOa2gQ9Cmzjb45noEyntIpiZodOs+5kFq/z0jXgldC
Po3i0gbAoMEZUakPKtV+12yieDdkXFkonS4MTOQtap/WFePkCAuxNmuDTfgjrvkSvmH8jtMU6IiA
am+3rUGc/OpSoohFCoSjTxMcW77wkEQ1CIShgIaHQzLwXJImy+Ce2yiwemnayK5Vgv1HI4iv1K4k
4xylK0eNTAkMoIlIKfjLF98/D6BnXn7ebGg0PTuHWq5XJTsoyEtZ3Jo3MC9oXa2V6Qoawanko7zC
benlobhtCYqJIyBjPUB/1vKgpE5OHr73cJhtCJptXmIHYaToETz1a2KHATji7ulpHjswZmd/8C44
4Uhi5RbyIRjYmspC5iYm+tx83BgZuCM/tAxGVY0PXsGIBaA2N9lThpMIjtMg1OYo3+Wk8qgQfPO9
afoetWIF8GA/5zrnq0RfVSKGjM+6SHUsuo1sXncnYCIX/27ejME760V608D6WnEZV+rfB/NsXzhu
2CI5jCfWy+vCbmI+3dlKomh5RUishFYstBGY+TEvV4QFBzmW82zuoXbayPVK5RpDK0y+2mccSA+n
vF192QA9yr5O/tHzDMNtPpdkVp8n+aamN9Q7/c2gcJuzCmB395khiRFzpDGAEre78PQqwj2lYCgQ
Cx5sSGaAFWgnITwTOT6STofKoZqhKwVRr848eNwrOFP5/WkTC7r/rEcSs7/S1X+bRIsp/emLGzgi
iA5tHKQgg2Iv1BK8iAULIEC/MeXywI3eaIYvg7d3RWZTl0JKWNBF8R7OXt/ha17fxKxPDFNRwjVI
NFoatEN5k8s9gmnq3KNhXjPpzl422uZKnsaOs5KjZo/+ILnZFG0KksafGpLGNa1fInjPhaxIryeB
mU/L5SP1sr/fxR5mIQGlWSeWxtcbd5HXx2xBrKaa66mdTZj/ARvWORoUG+HDY+oxZv8dh7UmyFTL
oQRXOv4nZxfvBCjLmPAVF74HmbG5W6Rl4sZ0YBZKp3HYdVCLsZ0uUKaXy52oCK2J57uE4tCFyjk3
fNJftQNtVOW7gbeD9Xgc0i0xd8Z3yo0OKCG4B2i/v9ceYdbU1gOog5p2q6KopwBjGNKnw3mDurfv
KI6YXwpn/LnixP2BTNF62vSlWuPHQX2aK4Gki6U51qZYcph8vuYkVqc6c0BYk81XUak+c663FFfc
ZuvcqfrwdQ0NnwTJf4167LoQXbV7JdgdSKid/Hcqx4QigBzpxI4E1GWJzOGbG2bQEayu++8m8a8y
Rc0SykX/9XaJeMfnzv39m+2PAcx6FJLspcq14WF8guqrZyBVxZ0x2ppXTfSAj5B4hwdGn6m8Upu2
wSv7okrI/gboEY/X1IiJarf/oX3IlUUCBXlgoQ6j1WZyfG41CLBiqKTwXgl9qUPK9L7E7ImT1wz0
zHx1yoLunrgskC0f7SyCU0PPwJuPEd/lDAkbPjzBI+HlUc7jOrd2IvycMgwf63cu5KXBQXuWftYV
WL5xERvZrVezgfHdJ+mYVVb8w5k5oGORlV8jXsPM8RT/MxhjOAr/0r5JWxDopW1AaC4ojlJLdCCK
AK94xpyWclpQxKF5IwPMaeJ24TSs3bQqlt4j5QlxOlejkw67Ch3EeMRl/gut13E7n+j/KhxUrFCo
ZIDCcbV1JiqioSv2C45+AphiL7BsTG+qBsyF6iInLPg4FnU5ILqZKSCpQcZbJqs5s/39VZgKRpkC
S0IzmezTnF1UXG8xkfaVGZsIXzxfCqVeb2jobqAJ/q3G/Nmvlo4X2lS49QPF3ujERpc6tluNjuHQ
p85wGkN2eOi6qKagSJcsJMSAP7J3cXeNmJJ2IzC8bQjzFsFZpIH+/Itg58xQbkIAXXOm6sj2lj3u
QfVGBCsznrLeRV3XYb18d/GSarOY5dXlNSVM+NiylZuj1NCMReUEhH77vj12iDKKdjk9rJcOSg6w
vpDSneC6qJMyo6up1cG+aUo5DhsY2qMtxiKKB8imD98cav1A7X2+Ql2SeEMKd/4Xajw/+WiQdfGP
WCDJzY6h0HbkG0dk3LUDeooBpZnmMNMwMRzNVqWb6ZYJYPNoXSqhtC77sT1Z2T2k/P98awPZ3qCw
JUShqbKVDpyaUzFJC8672uqXVQKtAHFLdlUfDa/YIneonoZ6A2+BkKdNgltqhc52aHo0XfHDdlYP
XWTNJQc0w6VqEx5Mt09+7KA5wtY/4u4urM2zY7g+Ay1srgVEabxdwyzlb/0lQjlrhmQS8+hSSQpy
7hD87aTJIPI5+EwcIV570YV5b1JYPge+ROhTIoKw37ptah5aOcrWBPiB8Sq02M/X7LtNLUKONyBn
RzDRr8UytG1YDczf1M0RrV89WvT971QSOjYIl6LYwglqbwtUyyheugSzVqL+XUymfXQ7bF2ILeVX
OshgRWn5Lyh6if3VmjlYlvCLcrx2UtT2UJOnf8YmKWHcxAGk6hf6oxDU/DK+1BvqY+XeSNCZt6rp
RToNYsrZuT5fd/PCnJpx6O83HYbGY7qW8CG1G2gJFhMYo1io7W5CHZp7rNKF9vQ6FpQJ6vZkITDt
2gUID0bkuqbIKpY4WMSxctOriOaJUozy2fF7XTDA0BjCyt2Zb1nM0V/5b0BJJ2KmZhQ2t2IlfVG3
wxbQdNchaS8Qpiu9tV9iITKXd+gB5cJSNM01l8GeuDbvw+v1abG8bOjCy63mmaDJUQioGzcrChuo
VI6HIdMlbAUIJ3Hdll99zE8X9iK1JsZ0DSHz/bIaddvybgVTZf/m5gFO2KojL8v4g2QXOt+pqSyK
jSTyHbWI03FNOKwDaqfxjuznVgXSlGpHemhze4p3/8XmucdYgd7gSsrT6OJ8lOMy8C5l2YgimY/t
9a9AWp+uL3Uoypxpx0lbK33debp42pZWxCLHGqu2eeuuYYdXneth88oOXrBSrUwYO4W1yvkQZVYf
30Gp5BlHdndrdrsWHE3loqarDf/w494YdMZK6O7cKNCNyQJVEcvDrPUSCYH47A6M5ONTnAOPXUaz
yryKJyn30uGk9OX8egmc+aMzFMoq6b1LAUN2q/wp2ojwDykVEp7smFpg1JSa/fjv7zPr/NEETsaC
6py3RP137Zb5klObfQy/KReuROuJisv9FfzdfJVnTwPGH1O2rVLDrUdOYIdVF+3ggQpWw2BOEY0H
fYvoyk3wfmeWiXrcdQIxlXLcDKsW/MGGHokBZ95R1Skv3DYDi+22XziYpEfy0zHQ1hz9m3g/k0Mr
HOjv/YnMS/t9uPdGkBy/qU5AQbmTYahGX5EjUizUYQErLWjHQQsdWrhewOKHUBMy5hpJE/zyfcqL
71k8IuX/nlHomA18aTORhQm6cyreDLq3z98KnKtwVx3z45AR9YA7uY+8mqsX7sdU0RvqihP/V9q5
CnpDnWmrm+YTMkZ+zjDMgVXmLflOvL06l0hu4o4+KHP8lwdMjrHUKQDw/94JdkLw2C+kX46O0slJ
nmjarAUUcbXYsHNh2aq2sXMvo3AcmBDrshfBuaQv3QQeRWhqcSuLvVSt7O1F9X0Lsfle/HoNP9Z6
7ndpY4u8UwD/TDM2wigJQiv2c+rMclH+f7QI9lNEIiLJlC7GJl9EC6KkbEQ2jqOdBRUa7P2v31Au
ZO2Q2lJtz3BhTib9s/tU1HrZKP8O3GSXKRDHJejV9uk8PlyXqko9zeFAuMLvei/nxtfydd9GDvcj
MeUxJ1PWNR49UKbg3DCi6zMEdKUyh/MSO5yylgfvlBy3LsAdQmE4cEajh8xq1Aq0B7EuNhzJbvdu
lRQgWuNapugFR7TLacOoIf11g3F2KNAUf1ge6eOwYTrSmuxcwfpeHwqOgnI7lvbOyFFYM1yTpWzq
v2FawS+PIPy7YhJ7KOHA7FBwp6aykU4feC1Qd0wkw0zLbS/nOy5LBXCJ4Yr3rIvnXwy7+OH3oGDi
K0bNFxKS+tu8EJ2yqnNj79CPKaXc6JSYuxHjo1vAGiZibVT4E2abId453b5Mdk09x8u9rCSAZckz
MI2aSzPxuHTLaZrIL5/ez+0KFI6kxP1XB+Coyyu1nccEQ51vjgBWbo2IA0zCUwmmx10XArcGkEC6
o38NeO33/ugd3buNHYJ6ZYvt6yd4OKR0cfopfJCPwojvV5ze+oJy3/7AE073c8z5vOqxLscz5diM
nKQXd22FWubujBQrYre2bzvXZwMpUfOZZ8lST3X4Bn6MZnvnAKnakRXrSABGzote87g0vVrQJeAp
61cQ0ZsYY9BGug9cOtDaM3hVxIM6M45vvUpRgQXo4598hDhlwZnzzHQ93mXwlJvON/o+fNeB7DiB
dfA23kYpf83Y5GEiBO6knGrk17SF34h/zH+Oy/wb9049GxysiJnQS6LYuLzUG8lT6Y0YHv1k2gH2
bdqpKB87K2L/MjoyUM5pmDu16/jy9vAfPr9giC+FORQ0NrgBM1wXkFAFfpW0XyCG0Jq/IZ4XJbW8
SdYY0bEv1rAJsL/686Mz05N92Oupr1PF8F/Q/Jw9k4/7Sb24HNaHTC3qF01x+vldyE/NSags82Uc
SRAH4DYoVL5kw3gDZKy4rvR4vS4dA66SQ2Qq/haqqK3AINPWyXWRfEPmpYWhqFzkQJiqWqGLV32+
9CR9QsJYUYpPZrcHXYFVHetsN9Vor8a7e2mYv4DYgpZQikzqAZuYbrq8/TnhTJWqA14OHy25vns1
Js59eeE/9AVTWIyUDYw8tuf1eu1IUSv/Z/aGtMFoBt5gzyqnaeDGU6cCWWNkeG80RpMlYFLFhoJ2
Bt+dNUt52E5wNUWZJJcmv/rBhyttJIkJq+RO5wgn1OMwoJwQDunpyaYK5cmDVzsLXd7paes22hWj
z7cwxQaGYVAlejUSI+TcR89OO6hzJmPaE3L5HIh8kE3n82p2pE0Er901N04dNK6dlAYPEMbGysQ+
+T+fAsHmWsfQSyl5FDYNjveyvlbvRV4lkpZLnFjyxF33Y1dYf7m9GXthr9s/7W604vwdMVk5g1tU
dmEG5huezN9zmMh3b3eyqX/c1MkT8gCiO9mKHd3pws3Sm4xke+kyJ5LasreAVUDMRSWqUiwMg+sG
3M2FTrICi6JHn2KfWiPHWS2u3QdOWIr62BD58ZPpOWYSUxv7wH7i3ElwCLqwa6Q4WEpJ2pUTxQ1t
eQgrYXG5LgeX5GGiDLJxvqUfYQwS0nNh4L7yamT6TMzFSX+295WYMA6d86S1T83kUZ8OtxysCMWY
178JPT3QaK+jaGz48Mz/fGrsTiAqlVki32UbMPmQyCj/3oiLU8tIix9l1YPEaBdcVqpQ3W/+dbxp
z0x3ufokDlxwj96R8Gd1/rzYEPq8RpAbv5dxSps+W84IBcLHYxUde+j2d+5KZ/s1B95lp5pga1jS
lCreND9iLkVhBI8Lo5wpKZ5nU+ir4EBYICsqZZZTKE8Kh9rPhMcFWTrphh1nKffB4IjrX9A8QJD2
TfUKBoA/mflAWDmMtkCP4mMDBHRVzr/Bu2HZk8ClFfc441rK8rqG7mfvPdfQCGFBW+a5OOWsIIjv
HJ3cDgypZOkmQ8OskU0Qml5+nuHdTVWJuy+/pQGLkElI3UUPTn3NjfxylOgTTkb1tyHKsfSOl25x
SFnlKbGLPU1vOyagGPxjkAMRVYq3Qm8IfoE9OViqZ7PeMYu4zGrNPo5QOSt0VwanXq990wOdOi82
4i3Cgs8Cg0XVUN5Wfp3fHkDRvUiKVU1g/hARPJnehfESh7P3VetpNM/Z3oiLHzrshIw3Ed5MY88p
XtrG2LciJlva1U2ju4Yxegz9wQy24p7SIvAutdVPAYp329qb57X/URjg8KXbeSDm4OaWdCaFKxsZ
ni16SsrS8beHg8HfLj+BmtOy/J5ah44xqC6fJAc32/yWP/z/MHary6SkVpXaClJSj5tY2widA3q0
DGSh/t/UOvlv/lFR0j50DpkBP5Zq5YjFSBgyBgGdmya/3c8B138zRGpGiWFdvBIujzyGm00M+kuu
RDnodH2fdWRWzscVf4ikxjfrbijO+vPejKd0o04HImdSdTuKsI1azg3EEsCU+SOEd0WqP6pMqIlq
02SDloroa2NgNn1xlq4ap2ND52kBsRzFe/B7IV2fLH1xg3rCoxhT2Se8cAknGb8ty0PSbW5zTDQf
OEtGsZqngDI4cjsCiYFFGjebWnv6+j2SS3M3jid4Bb2a+Z/hL6R+3cY86AS9ZK/CSEr//N63N4Jk
wCbJO0KwB4ccjuCoPO+/DF5OiKIGjAA8toruEZVg7DKT0LMtK64uTCCTIGlyI3pWfPQxG6FkPFUa
MMaFRu3MRFi/sBmulGdhUyJ9yj6OjI+k8XbE7vtvpM0qz+XH4zf+1Eqj9AnOEtqJI/bA1iz5rHv2
QXSbRiRl7XPWHO6aaIypVRQglG2VkptCoayKOryPhJFXIJSqi+6CpyKHT6WHmo1yKFx3GEI2X64t
ibX9aXB1D0lsvYvtYTYfEmIEWMnOcDjdHGSO61rN5X2PFI+x2d0n0xWga1B58VvTVps2kfxCaD9i
YO0YqEYoCv0Q3PjYSzI7TIAdbmnNdzr9m43anj6K9U3J35XWyfB1Gek97LlfGVxszsrkRxsrtCHp
rcdZoCD7LWBQz6pUUrglqh3yF9uJxfPirAmxPwaUoKNvIIELa2jS6dATTsvI1X8NJklnBiorcY0H
NOP+Zb2XEYIwI+aEeADe94OTg4HVN9txchJtg2v5PYahM+Uyu5t6odXBhHCkOya7bkmEUPTuz/zs
d5lx6vdwE0jR8wLisTpUWPjSfSEKti/IgK3Fn66oVeG5ct5A+Dfx23l4hVo8ac2PucENqOlZccJA
YV98HNFVELjgm+OTzSuU2Aj0e6SuNcuXqhWSMaVojcOWcOusFJZxxCAz3kleX1GOc9uRS9iCECQd
A7IvXJFgjRqHW1jt2oXyiNF98Ngc2ah2gW8c2X33H3ApGi2WW4SFVybG5ELLoeqerFq2nHSU21Xj
9esmo/HOfMyIa+LZ+gulespL0O2pCe2wnHBIKoTQPSvBxP8jJkNgkWRMvmV2txQejDWQhimpDKre
CM2+yTp1+qTtcIr9Xu2XLIUJt8ve3JPiIQTI6QuVseYCjdcVAuvOGqUctoUZcNrY3VJjaaNoFy/+
SHMPdYJ+NHePl4fcucK9LKBWhHmQOSZsePC7qohJA+0JiwxDHKMu1AyVjUgHiUE2oI0AuZ+xCtwO
0W2GuAUnv/ls44CMYOyXJ6AO4B3mmYJ6hs+Ry5Q0/imC1mPaO6nUDZOC55fb/PlFh/uKG0ej0f12
x9Nia9RioGx2UvjffMX3ErEzg+/UvI2wL1l3lkh8qfk2YlbKCNAj+fEa4mFAQb4pUOXBQde+xFDX
qjk1hNarCBjaDoP5yhuRE2jHYv+uThVEITrnUhSujdEAa/J93dad1T1aK9biEeEK1ToIvIObM4Th
lGZq+77Djn+/Tr/NvzMGtebqw5Um2G3IysFtfNg8y/6TYfIi5cQuJz1Ed7nniifPTtnQObEvwoct
RZiInLy+6blXS8D0r+Jso1tR/hlnPSR/Zx+bi16en4Ikj8/vcoC3Yusn1ggaqXub0+PRdYgCZP/2
76p6jpdOsAX+P9DORUz/h2Gk5n31pJjU8vGpVLmf1KRHX4XQ7RMjoxw5tu6wp53HgJXSrPQX8ZDo
UmwsbfCB1t5WAWHPzM37mLOH7wBwqb4t6Dw74+gJcV7BzWK4EtnuAOQ7dr8iU2IfsVrQPkzV9GDe
iu6SKydAExj828Km75jgNo2RcqZQffG/X+gIi/z9UU/LTr0ge9AWeNmnWyf5WOks3hEJ3shDYo4D
9YJucrFoggeMIeV1cgVzpzHKgLZoUq3uB3XmEj9DT5VPfR2EzGJzfJhM5z+1lRN7Dm2hgK6FRD5p
oZvj0bbESdiixcw5aFfSFWoRVueWu0PVTGYhg+bJisLsNto5AQAVmC38msqgTiRm+DsAFbOwXeMb
Pf1vqhmTfz74D42Pc2s4xQ1bAgmkFiUObGhuvyQ5Tw5kpOjDXpp6VdmCCqy53/X6Ej+feVkxL3W2
Zf2nIP97CmU35vSzLQNSDQ4Too6KBlxmV9cwnNxNld8544uDuUZHucHpfKj2yVkB8CszF6Ftxl+h
Hd+HFi/VFcCoxDJQkQrIWoorfVkCLCupOJNVYgUcZszg41QwoYsaGVACPF496A+Uxz5F+vEsCGI1
lG7qBEG8PK+QPajAS0MrARHMeYGg0OZIKlQwHVxYqQIm6/tAZ6+Cp95fZKegtSDn4f3Q4FFa0lE1
0NtRUAxbimXQh22D5p2DS+uNV87i0nXWBvhPBqc1DQNVmp9Xu7LcSDZD8RKZP7iRad7Z7tjAoa3c
TTnP4OSEz5fSl4vlP4B9VX/XISaB5SUO9MF0DikTCR+N0gAdxIbf3RWvU702mtIsD+EoFD+5ZU25
M9tZsIciZxZELELIgkJk01ozVc2M7JWDw+8D01EFI+6eypBf/9bJC2b2Q6srP1FWE1n1EIMPtvhn
ZyNipb1knnfik4oqoeHybra2Go8PjsEKPO6m1NcKFCj8FUvGCzwK5kPeFzZNfHybf3VlZetpM3Sh
edeqv9VuJsTBE/TovP43sqwKi3XMhbnbae9uCCLJR0Noz5ubKmQfWDSS9h3jxFrehO6F1G9Xz7FH
jESHkH5EFwQ789c01XXSjf3mjELo2HjWh+VLXegZEgjXTcu5/yL0eNyM/0sG8FZnSaM6U0JJFwBg
pBFHmkjB9UjtbN6P+TMf4NNoegGpDhgKDF6IgJ6K3UgUSokFJeymc+9qISF5AdEGro1qA+Q8FXt1
8T3OCbmbwn8PxuHgrCenQmnSUoEShzwRVSccOj6sptLZNEzVLV77JIxDYaZaOBrNdt0WLsRM3JIR
0+2K+wp0S0glG9ksU3IXLUlcFjnxpccgWLSjqGeLlq7nORgQYCBZYwp4v4a3lkUvD1fQeuJDJ1Pt
XHgTjaJc/9CoGoUb2R0dJDjo07NnolK4jpLj9PTXsK75CYrh0n4SZ1MYK1BTmDSld9BEAntwr0P9
eS1pXFQor0FF+uWgd5MA8vOAAP4XRrMo1zdrdZHGrTjqBW0mjDSEQUERThWDPbGvCg88lVmLfkPY
8eWFId/+CvvTQI6EMrWbLtxDIkrW/ADDiq08FdACTHKHe7IPpLC/rarIZYcglRiwniuOcqhjDPZt
eOJk1uj7aS8uvFgmlVR9JvjZV1b4v1CVN7+3dhRxsCIaIPW5iJXCOHRcI68rGC4/Ljxb4MMZ/l3o
HsUgQX+aCFIqxWtLxxDzK3c5or8fP4gM6GsczRkZVZBt+9z44ju1cN2MxJpNJF9aJjJTaNNaVCWZ
ssS8BtjQr9/sg/j/30E22Npd309nwSFOZbgl+oIvhl2mvpCYSBfP26wbAUI3al4i1f0tdRRJVJts
PWgFonV9BDhURM0n9+4G4f25J1wb0eNB5VK1xPyNNX9yEE2SVHGRBjHozxTF19+nWyWc7N/lIUCx
02K26t2AB6faxolKFlYJcNKtXUucjCD2ROZ6fkuLvKtdY5+l+4aToUANE50XFaA5pwexdwUfOFAe
otr0pV94nGtvytrLZOB5bA1QnqalQ7GlDtAa3oVZCljWMslb135xNdePh7Xuo2EvJOHzD4cVoeFM
DnyUsVheYLNIaPveVCnAqOAaI872xeGXkaVRl06/5MbmpOXNFOOn5Nv+2yJvDnu6+JrOEOwOwPIt
fypEbPghruh9PdnnQY0VhGC0d5HSeNv3CKwg0YBg+7l2/ZRiJMqwW7UmxDh1SQGxpj+SNxhAhwYw
OEEbtI3AJVzpsjj2zhCxp5BSMVgP8UTlskAMcZ5emxYJ428Cxb0wKPh1jLPVJbP8VU0z4F7F2OdW
9SUP5pcCdOm/2VSfNMdHmuDF4i92flOKXyAgPV8+rVakqyJ+FYlKhQse8ac3r8JjMHaEkiF59hRY
aMDdADG0zktQ43O6rcjXFWVO05SQVsq5CAByeKA4wiNB3K63Cna22Q3MtHxi0kj9Ct1maOWjaUOA
6AZDgxObgGajKcYzoWoULH4uv0WjzTdsaSZFDyxWUNP+jf46B4b5tVakC/U0Npdw7tXN3FiuKVnq
DLkXHyhOAEQSvxjmtS3U1MFbmwcBYlV8tG4C9Zj6QhE4jXtm1wf2fB4GtuRljysfxTgXdP0VOUtu
qUzNIjAynAHBruBZzKgukMdqJpMkhYvd0gh9MguhXPd5Q2wkLQuR5JLPRiEDGWW8Blu/XXQw/jie
eCwJWRcQ/lNa3ua2d0gWyPVYz8vENxdY0tbGEjYphya4Z87D7ua3iZ9zjtRR5EtzbAoPM7q2pqMO
rr+Lu9dxzN3e5ExVRE4StS7mGznPb6nfmi+VmQoAaZX2h+l1lToS779Fm4XXEhA2QWodsE+7jQPb
IkfA4WH4jS6dEkdDCwImyO/0mn8muQjOfVR0NBt+bVU7pg7gulv4UNgFQZaP6JSv9oQEa35ndwSz
Yi8fCNmaD/Lf3S3AyLAIH3B4XU16ssuNmgxgwVz3PFXjZ7fNgc2RFXe+pvYzVRPb5VA405LaaY1L
rE+yUjpTpeR355HXrldg+3plIYa3e7XGVaphXzwyvqUjJPCkdd8KbjL0Rp3Jkf+KfDMUx4/XLYp9
LUw1S7hoBarsSsE1YvKfjPQ/3rZOLX67VX3PlkeIg02Y42Eez8L3zC95AM8RMhSK0voy2nz0/53b
R2RT46SYJLsTaOwD5qZ45m1XHlNqITIZr62Jo9o7dQINlyIY22Y89TplPgpqu/K48IGgnDlHQuN3
yYPg/01cHfUyqYg1aeE80tpXnuxBXXbiEi9hP7w1Rs13z8t/4KxBuMu0Ic0OFZEWOH2lfpm1PMSS
yMNsCbacz/Mz/m7SnunkrRF55SWky1ihBHod38AOL7lVpBm83bwxcfqMM0Re7O1St/KgrwhY+mxc
t7r2vFldtuugpyqxyGn2o57HRUUWaCJ3AS28OfjbjPSC1fB83UHzX3HADhqGNYqcmjYV9XurYeA+
uW9t3ZtWeySxe14UucWOvKVGlyZuDdSGYnh0kZhwrrQeFy0FVBZIvhJ0gDJAetkd6f+Ne5wQXIuG
JaVYkBqG2u4a8UCBDjAnSUetXXfhH9L9/5Xs3sSk+gUSvTJPupyh3mttAYnPFFExNcY+LqaicUL+
JCOEtvu3sNtL6jk9Gjqak9fZTzoUJ0enPi/6Jh37Vnmw1rd8UQZ+J8CAoZjDwI+wMrNDbYWmKBcL
MEJtEsdbW9jbZRlgEJJnUtROHad6MiZ3OAEaRwDY5evWovXD/Zg03+1z9EI0a3cYTHjLkSFp59VI
LJlnGuTFuBIxhGVBzJLfd/D99b0ZAtOcqX2jvt+O04iSVNcSGbEt0KZp36oy4GtrK+NCaPfQbttC
2XuuTkTDp1sa6Tm6yA7ldgwODSf1HlUTIQy7L/w3C7y5uwhT4VAn6s50uqayZJTGUzE9TZSfNAcS
rr8mVT74h5j6BUyKPbPzsqefqv6P4jtLMIhiOyjKTdQz9JwPoIFulSY++3oWqIu2kESeISf6+Pok
wZg27pMIFtn+0vxRiKbaNnbjg4Cu1CXVfzTL3Nve6Q6SZXphnOZwyxMEOW4frkm24I5yCnghqDEF
VibLb9JsvDUAKkB0tEprKMmN2URo7aJXAaelTLuJ0lgORZgbd6Ud/WKptL8jLv/hVVaJ7shwtg+E
ZUmSkmxJbNxcFTKVAppnRK105GQHFTHyNleSmtOboGy7RxZzDUN6kprzn6GjwcrAzSqhxcl3N0KD
HxjV1CaHhM8b0W3kFNQHprkgWaZZNsgRXXIeDZXnZQ4DOzP54QJUQV648jMvw//zlCU1eFst3OCi
2jsXPVxwfJzjncCLjja8LWvZrQ/h2IVRmmwJ2pnu/rvOkeEKcP/wyt1V8l2Y0e5lkbQvBKQqO8nw
dUg9J0y1rN+Jt+POAug4ZPHiYAoiN86IjoKCTxgGuB/kMAAoRawgYwgxJbYNZ2UQHPdHbC28uWVP
tuOvNryOQJXEQBelbAomsk4QK7bjPgxkH8dc/fq5KpLbYY3iYCoL3+jZlupbTsNbw+sdutmSBPES
s94n+U3lJX/36Z7Yf2Zo4hpGbitNpfLBGmQimtGIxKiDKKURQHUqRmSYFsWX/XsQnTukV/92/5Vo
2DL2sWZq8wGkjGLtMbaMbcatXOWKMBZBWpDYlK5up8C884vKsql5HfmlsiJmQ1P8W7FLF5B2coBP
oc03HdxDTUg8r+vD9KGGu7m/aKJiPkoKmW2MXPYc8qbDeOohwIIpzt0WY54CoWpojrzJAop4kIaA
3jwuL23+9ZKylWw16lMpX4Pgzt23DFRR+FiPyftD085l13lGq2gwcGcmM/7vkjRMIe4yFlKWmyLp
vra05tEIS0XkqvexCfxTwdf7/euQjaFTSHeff73XDnyLoiMuVOKavbE1/9c0GOzFFeT6C0gcPeuT
moB2muo4imOMX7PvxLWNAKrQKuFDh8AGEgDa4Jipo8mfSOAg4GHu5USMJWQQCvVFRUT04+8XH+EZ
tk7FSbXDb+xxVpxa0QGE4OSff4CvTzlSmJC1NUuaF0cjsoOZVQp6SoPDEAU6DcA0TpdYF3iUuERb
LTH1PmPZcf/8WqDdN3e43h4L4KINTsiAIXtc67pWNPiItFwlw9RZDghRmP7L/JV3m6Qksn6ZigWg
VH65eRC6WQzozR4CAWF+53DfSFH1H7hAIDo44fTsHt/BSTKdKmX8CBsf116FfssMPB+zf8kfgozx
IOTkScmu3jAYPuPVZxjIVaPTsKNmNYfz8/RtXIw34Z0ujWDPk8OE/3Q6ZZbFQQkcsmrsYWvetmoi
60MRVI99hGhFWjgvBX1beO+gr2E3mFBlS5C5CtPOjdIvTt5KOL4xERhKcVe189oaPWJ2rbdUwX1C
VnYzlTx0f3flPkFT1vmJw3uYP6h6e7FKwaaq4X770YV6KbgbRCbmBHS6wnbFUTA38rgav1bXjruE
9CaFg3PwkrsCXeZ/5YkGQBqnmBtBtNFrvO4UB++XRBdMfK4PuJbYcVb0TQ8Fh6t93fQatZOrQbNq
cGlUBD5uPjpUFYAUOZHavSKSPaard7KFFaDhK1gn99NfvKKllxQfOs5+nvFXbijkd4+GisLhQuDu
YZOY1WlHMuWE96frMovU+cu6vdnB3y5DcuAB56I5OTMD83kk7/DQI9FLDO4kcPluL49rBgzYmsI8
IWIdUAsSuPaYHmBvH7ID+mpJ3aBvuoopTVXvh738pmoXMvxVL+uAwE8PL5IKaIdeEyw1qN53RqvT
RkVSfjo8dQ4FJ37lo3VMgAdRtirgn+pjNCX95+WERt9OBImnmUTwd0MVckQeZHj+SqjdXGUXMgKJ
6n/s2ENGoFZmLAYK/IcMcgofVzr7LkccyJyVRjrcK3uvWfMx4OAEsQOXE6gmxJpzVLc2SsmcAo0X
n+YHTfB8ry+oRRcN80Rn9FzPFykoKWthS9RrcMdceKC1fFjtgEQYFA28LxS7Tfvij9MURyrd/Ffo
E2svvgSWdf9hX2ARQEc2paiFUeK1XcId+tL6xWOji3Lunlp88QESsdJ+gQOsCfM7ooEj5tMP57Gl
jr/pVPmPpzXOR0pqdzLkllGt+rJJxQa4UHNlCAdNSZPGljXFJB0955HE3AXwtFS3kt1v4Y0587tc
FtPTFVP/TUqltlp6yZ+B3WrgUG6NYnUVgQNmOJHixVPrUEJOUkDXNrbWpJW6uk6qaO5dgwhoQd5m
VTEk//eDOv0xCxysqT8/ffYvCxlTD2BNdc1pv67oVJh77RUmpOnegZC8u27C/iNN9Hf8epZ1673E
9zntHwVn9oXYiKwrCEzWtQqmJ6WzoRnnGz79na5m+WKNyY56/IupjFl/FnBNRQUmk9GKOaGpnE7Q
3Mlmy0+BZAZ8e4CATJY1FR2vQ/IQJsZvWiz4LkxQfIj/j3dIk0ezI6S6ZEa9rhYX8JMhTl9eccXF
LbVdQwt9Kmw3mEpS/kiVVKoOhG1N80Qs0Ne/U1+PMfQWVYMmjjdiD1iSExCGdSL1G2b/KY6LjQZ8
Q3f4UExUdW3+RJ5zyTo4YMvbwiPzveufU7Jf2u9he6NxYxZLJQLxcHSCjRfiCtZOtqpWkLL9A6/7
+bmyDSwAOeKcncGtKUNV0jVWdYZNk017NeTD+PVWDqPNS0eFBoSdP2Peox4CPjdfCUs3dbLqXBlM
r055YYd3sMHx2y70yN80+3XfF4YtQUgd2Sq+V0fjsko/MrZsrlb6UOFT/J63Y3wv8TQ7oP4OIHai
aBqLTCeHeEU6AnBXJzpMPse8GHcj5OjqZmHjIIUcdSFFt9PU9xry99vPaMjnVjpwG0C6lPo/+9nd
wiN0uy/4HtgvOUzUMHCU4gPZFTzcvr62sV6PCkLezpcwKxrHFX4UXif9coTkRWTbRQq445mXrIeK
JQeg7aHstFSdps4L2+Wakk1nsbeYfe48FlWXGwG1EAqrsO3nks+8TiHnkCLrlOuLfKUFn201kX83
JvrSUa38cpx/mtdSikEN7dTQ+WWxjAzm3BzstNlr9aZHSHXqn5zpBitn+WrG+2oj6vbXajBai9sC
wUk01I3bgyo/MFwrekKaZL7Do8c/tes5EHJp6NMm8oaKSHRJn3ThxAXNdzxR6XDwSaw3T0BycohV
Ysu0HkQNI4JPwciEdmkbWRrVg0cd6LB69Z5Az+Av6jffNB2PQoQJw7aLIIbcVYizUoYyGqL/q/c6
evNKl3tJCot0qhleFKzsaukvRx7ByiV2aUliSKWGyICMNejWD8DgWUi9EF8c4iTbm0n9RcNVwQrQ
CkzpEjtHpnpOovAAx22BiIVWpOmsJOjqryKOYYuAQa3vOMEuJq8XElur5UulvCJ3btZVniykK0Cw
Kqryg4PMkFYuPws60DUd9roahfNOqEqMx0UGUmb4du8PctorYz7qAIk3bseORxWtfTpg9cUa1dnZ
bKeWeJwV5ypr2mDo/6Uo1Xj5+DlTpqACdH105/GFD4mW76z9mA7zUT0EUFee8HsnjcNFAbwmVZ6D
O+qaWe92QMkP9hbCMDVcodJKXwefGpNVsu79sryfZxQrcBE1EMrfBrHUBKskOuaqz0uLk6AhamGO
y+upKKeryCIL7di7JJGZwi7JXuu0qVTK/pAjXVLa3RkaXVVX+HQMEyFSkLkUQKTEz5UlyN4O9Fma
Ba1nsToO8znDKxULDJMfBszH+gzZ/Dc6LMXot8zlnJvBV6hMbXxJrDzqOBXAnR3h0+shq/aaGnU+
OwZzrt5VygihB6PrcuenkpcdIcysXOitDRqMYDKkdv5OKM7tCG3vZ+vpo1OXs7R1mYoGq/PcHaPy
+JVtrwfztfokR7gfjTyn1cCeDCmUaS/qOZcXV7F9U4PKtsUyRUocf+4cUBFwvtQIPPnspAMGwCEy
hD5Ufrim2WrHQvkefrsWyHxghp2BLFIXZAnGmqu0u/xBuPnzS0PKXEXW6IMJsFjWI80mAaZTvut/
5cFdNxUm1Q4vVbTX2mHJJ7fkC01TR1YoNsH2MGxTdZ8MCkJxCBmMAYc7XV3mYW913WJkCupMx2BZ
55bi9onABVBcIJ8dKPGGxdSQ0iYqsvwKrGpIMAXRP7cdI3kdCF5pwUWr6iDNI5TQuIzjCeu3cL6R
H7Mz6FIWE3Wao5ZkHkJ/zGoxJ+pXGPhnycWQacxU1sQGiJLQeiU2uXWoFnhOKa6D6+zYJW7CFBnq
RhiyaIz2Uk+25uRiVGyHpoK5aV8oq6HeK43BIJDWkIWMXbKtRzKf6iLiY1DtxDXZKrrto10s/7qQ
8e42PEJaVZJOTzP5f0fh91R2yvjYuAa9VwN7VF+Xk8N4S7IJ68KWqZZJqqBleagkiYsB+NP3Dk2x
jjojsMu+Io+7uzGBESQ96KWjL8ZsuSyQtY+tkrOCU5H6plNdzB2fLuo792nlg0vmF4Fm79aQzgYk
e0q0dAuRy3kh3sq1+z66GdZhl8/YJc0YeqCUcwS8py7KElYMytBhtPJS90rvlR7alGCyhaWjEy9u
L/9sC6dZB1iOoEWp8Hntl5tus72zvueyUWXBo26U7Tm5zhiZ6qHZocTMBgZdKSK9nbBFY77CSy1F
yPX7tIb0vMcw3NvOE1BvX7caH6JQQ/jOdT3vjX9T3hrROmkDzCSnj+mt30umCr9f67wd4dz+MoQ7
ziibVLrgyQCnIF+ix7u18PTppon3bi7RJnqWJ88NxpncinXyvU7W9bvgRhaqYcMsd+NFfLt77FSQ
pKSfyXuxYeuXyJ6J5shmoftW/GM0cXxxXTwa1pgVu0r/gVKUhDx6Vci/f8QwwAJVhdP5oQEbAbdR
x3uNPUiAfxpWRjTexbd3ZIqfQVNWPqmVIIq3aKizKQaZKyGHQrdqfU273vJH9qS7R0EuITGrVDdd
l2AWrWqNqFoe2Jc3uwMd06mDFYNwJZyWQCOkAP32aoNMCaErco9vuy+WYpVc9rpijNw476XMFt25
61kJJofBMguok+WNZtVdWZ4RQK+vUIo0YkSWjZ1zuWU/EzeuWNzprBzEMuEbk1xry9Y0KXSdNivi
E0OGLg2yj7LeE+dxW93gMVp6wOmd5Rc9hUIuPBYdOr+ZEFJLTgbag4X5l8HZrd9doaZoQHPRurhe
dSYA6wEV7wNYqagRNx2UfgNzhnENmIw5DZYB8Rgr4g/uleJPSqUItFO1ZQfOzrkXPXk7UEro/Lx0
3HezOI8xHqVkWr+DuQwWfuzJYaoKnF4yfLee+v0zfPVSGTMjgeIOMOO/iKcjP7d+VO8ALYWD4sUE
5LvDXIwb8lupURL6v9+FieNEgmiljF502LuVO4/lUVYkm2HTa4ombMkHmUv8vkjsy/76k0si6pll
CtiSuudeijF8zOT559ayM+Er2uyvtO+ChleaiCyndYvAJq0TnEDteLW3T0b5HQKKppsI9RPOLo0G
G95I2WTZaFA21gxyxFNkg2qiqrDfC1V4p+wmF2hALOGRqcwLaaUxNue9bmg2SpLFIKU/99sQho+D
N4fRwFxWUnoeQq+ZT/7URT3qjDsI8VtrgCmZWdqoXkg9Z5AN32lHLaPUEbm5rNfK6m6vTX1r3osa
0muIxWa+UNEcCTIHtOGIMi+egI4iSF0U8aPBFxsEv+ZxoghoA44aeOA1BIDh9IgrjcpH1oP25Kpt
wMgFmfJbSb4wLCM95y7EJHITjC2X9Qpx/RP7Qu871D+OqnR9t38UHYReIG0HZ/VBOrVcRJ6Ji6kO
yInzQsyoP67daOjNaXHlxhBpzYuweCYtG47qrPu4cvCVAgALSrnYBr70re/m77yStUbfN3hl5k8G
mwZkYkT0kb0vVUfvAKjgpsv7EdiD3GOe0hYJS9O4DIpNESye/63SsGKEHyXi6Ot+9WSgXoi712wt
aLu5CFzTcg3duSgNiDCjOS59ZB0eUb1QGsB1YOW7TkT9BoIZvlqExYIDucBI2IkKtJEOFrklF+Un
qggW37u7DQe7pnVEIZYUX7wJR9TjIrecxcghye//28hCxCLRYyKj4zRMPi3rdy0YSfja4gRjn/gc
qEy6SlLZmlwZb2V4E1Y0GzRCdeZOxovK1w4CE9iBHFajNaoRSegAHonTUg27wU2/0YytwfRyXecr
IqXgcRcK3AvwURjaX8F1fr9+98mbESSd5bHOOIHiIBzqi5ITxqrOmmQL0UGlT2JoLC/guLQn5DGw
/X8R/KkMRypqhYZZZeiPFTTyyXgloErjgBx8iWPbock+IS5S0+IJc6dlnKazYuSRYKwEEHoLWc7Z
Cg0GQBZngOWVk37x53wZlP2KWv5JRGqZ2hWS6s9cVcZD0T7Ta00j90mzFkW4T0lAeyOH1Vyo/H63
gwrwWJsrXruGhskvM3c+wuIBdqMDJ0p7sRe8SZuVyB7nRtzFmrp/mOVYQj/gB9+RxWeH8Yovtg/W
StECgei2zOat69YTMyTYyTRWu1BtDhX7hbKGEgPvlymVwhYq3l4YV2EeBBLTokCK/IXdthefgOKO
xJpimvvkojO1o0gpQf9YaF1lOXMeYloJaCtN8M618Hn0T2IvOdgntFKp4/nUSlk5V8V8ArBnsila
duN2BH6sDx2WE01PJ/+vDeB8sM0zQUSi7gXXQyYCcquzeLSCyyoMFtPO+3rvIczzVoedMBpBM1D3
6jadIaQk4EsOP3eIxw/1uWN5HV5gLxHPfCEViMCIJh9HAMZIz/6yM26Jw9mHOmFMJF8HNYAGlYmm
0QlNwZ34SIMOf8usTG6v98Cxt50c9UjxaoO/BQOfItYiXHQrOZq8ydKIt6bJBqyqdgfIDGw977gx
UPTA1mz1GdNkxrX7VECVtopbj+L4t289B1ohzn3tTmdHyxDVXQMCZM2zL/spniUXZhiPCJZV+VUn
9oFKsyV1RzTwB/XKbqXW1YUohieU/bXVf/rKF7GEtMhtP4qm0LCjeU/WiCDHOmbafZrWDikvb1Uy
rkFIhdmmJxDgJ1ZzDCinsG+Jjnwb1+pGimFH8sNdaSqOwRUmD8Iycf8P0VkhHmFmnuFnnqJFPl2c
SAGkSuh9uuWKBQvdKEoD1lUfCpanw7ulI/9bXomf0yg+7GxnQStLgDzCvGWgH/i1PhtCkU4NX0qB
+tl26IJBHamlA9QgX0HVG9/aZhnhAzu++O42oANZL3k803O/ZYCy4m3D8qBJyF0BxTjM6rqzSWgr
7xRf3vca2jxlA1lFjtXVia395rWYpgfsbpHaxFtX20//z9aGYJuLyS8OSsnEOaoAnz1nw5gNTtvN
L2vzPtfZYkNpl64WKx2nxpP5demZ/ZXWhuDuhdhCVL5JgXg+TgeXZEJ12ywarI7CKNt6OuOvi45U
MFe5mJeZgIiqD3n6xI+3mx6ge6MQXrOyP1gKyWfGvzh1iFpH1fhdLufFJQHlwsuohdJ0AMn/+BuB
TrY8rL1JYxZXS11XoBaqJKJ9RxDLo8MpHItoQWwfSdl54iD8v2C9q01QM+2Af1+5XAoki3PCEYCG
vBnw+uajPCgMwVuJRp6+YaNTgbKwYD5uihYE9o6fUZSQlYoIm6fRqXVH0nYz/xIN6fUReHwSRo5j
I1L6IwMrD+YWKF/2jd2vSg52DF+uk4kLtftHVhhgAhEyUovxFi2KhUKaMh+/71E/fZ3OM0nXPFi3
KI7h4ZSXp5yNgGyWpsUesG1umEwcGEg3+aDAfzb2fU02zF43FQbeWUcfiiJSIhnjFWqfC0lvFStV
i+QWMpFPWjPaIAUaaM20jy5zsaujKjZAmWgShupLIakQTFGjElyTKaEL1hz46eEAdxlVb6/zwNet
DYRJmI5Nlgd4bj1cBtPM9y7STdMU6UvUUMxiG5hCPq4DuZ1qgucTeKnpgj2zQjnvAFUPzhKtEEpD
7Ym42HzQgC7KiOy/cP78dAYPotlh4/ntC8hfgadIARzumNxMljzWUqT9zUN1wv5BGZXrPj8dugrP
fzY5ZbHxeHBweAFEXeeQKTjpl7eGHXS/Wh+rRGZV4N8r6IFkXOWAPd7AsCwWernFDZOsy44yZq+p
a6G3+G++Tmic61yE5GLeVqHVtjeiT5x2Rev+NsR7hD+81hRnQ40zhJriv0BuHW8Ztkc6nIGv8c7G
9YP/qa67thOvC7ljobuc00RVnb6n6mBXdyD1AGL/zW22yBwi8Frni8S0cbE7Y7qjHk+rkfFg8rZF
YF9vo/oteSWsy6nnSth70FwQDzMYYRIAj0z4hWrZWPE/R2fmu7WWLTdYXeIoAa6ytMjxRBmLu4qe
H7fr9jwxvlbm/RObgHGUEQ8CeQzM7e880IWHrsw98ZGjuZnH7DBN9K3Ro8hW+QVWXa2cTsuGuYXk
VGJQLXsh53IqZMke1yhE4B8mtQhELn3UEDNRh0NlNLSB80enodVaaBWpl7GM10sEAN2vaXktdm9E
8rSmx8g6cPm+/MFtd8a7aEe9Yv5d9HX3+5q0aTNHw23RM+e4XP2nZGPOMZoFtM/7rxZSz5CBthhv
jyKV48FMaMdeqF85OMUxy70GNrVyvLBI6Kkh/A3QDbiu+wNr3eIawts1/QFX/OzXBfl8PnUzs24j
p676oMyzoAZ+gqZdUvwmuKd6bNayJ1Q6fqU5OU2WLGFKrMq4MfH9Pt+aJCA33qvWZ7m5jnhmnHbr
8oQgvZRdQ5xNNwefTVaD5/lFaEoP6r4tFZgcR/0snBVc1WYC4G+oULXVbxemsIIfpq1DoPAsJf01
GxO9ybeybE2Cr7/RZwfEkvbEddxElLdpSxhi+oi1HBnPCzqtyi6tCWQBsM0u0idzKdmWiDU8gqvx
38WliWnUbgGI6xuRp1QKdfi8FWV6l2y7XV6dPdpbfyGtKWSsepjgKR+P50M8+dvP6bOtQvyFFp0f
pWAC+OxYNMOrlwh2f7DgHhi5vfqK62cOrYoBQFJOQsNLMgxZBMyE9RcFnwRu3ELZbduWsUatXXMj
NNE49rUxx3T0JgkPfBjX5+pCN3v9TZLeOO4IXrsug/5MjYPPlZZteh2VCO7lFlbyps/cFOoqB8ZE
C3NKpJ+e/qZQwXKY0Y/o6hFumhlh9e/hDqLhQxBP83Y1deXFMXp8Zus1Xw8RGYiFm0PKHykP4f9S
y9m5RMA1D3CqFInX4iQXLgNuC2P4Z4xn1K/wtb6AUfq3brwLwQlcw9MsV4qFEtXeUrkeQptc+OG2
zc8uwge4RIBGef0RGZAUxXeX1rRUo+/YL8Q1lRDp7kULn7va2tB2FH+m3PbcidUul6hxKmC4Mswc
m7Jn0lOrDI/MtpdhBX41tB4/org6a+0qS+0Kol2cZbq2GkpoA79aaqi8Qu2bphB8wlsjuqhfkUD+
n7p1+x0TDSJvYFyFXulo28I1Z1hlx9kSsv3rxXWqJZI9hhDFVRNn6jwGJdJWo6LNgyIjfB90EIs+
dTR4B4dZy+Z9HzADHPHeDwpZEjJ/ZapqFbbTATvJPIbthOwjRQAVaqyp4ka+BvvbDG1CGJhYS7LO
1G9HJD0Obztoye1YGGx/HwqQ81N/QCn3yh9C+/HwOVI4Rg4V9vX2/xrehON+qHcx66MG9NNPtC3z
YVgLQ5NuPcACTuxOWi+VeUMi8ROSiflSddHXkI8Vxg372imi0eyQ3Xq7avJMBbM0izPloHdn6usO
wVfbodYVr4UgaxZIAXvER6cgPu9R9QGNqQPMvWHJM4AKswBZOz32bv7XbOPubVNlBWkLjYW1Dz/2
JSxOjddXx3/jxyLKZ6FnbIae1zWUdIrOhxeaygFx1SZgORM3iuJ+rqjZcpgzJzEe9/qvlbdEOt7A
hK4DuPzsiK3gjNJourfAI4wdrU0ZuJsr1cl3bPqaKe/1TFHcGWS1Gw0lvdtXwUgg3xZRnIj4BZF4
6UxxwE6gn61f5FkfI647HNfrOr+9L9FYHzJ1VmLteK6N/uz96aRw6mBvtMJMuPnluRl0b/xnpp2u
ffxHGehkySMyGPUcYXcWQW1BdfdO5uPmORvceZQUChgeE3/Wv1yCE4eTufmHwaY5qttPdRzkzExt
61ezKKa9FrAMbAMDH6e8IUDFQNjVCSKJmjJySHCPWMamnC8AYSzCu4hkGXxrUlyQ6EAmgCpWyPHp
HfY8iyANyFCt/MOY/lEr7CqNzcypA6d+eu+nJ6Pf5c7eTAZkicTfnO6IeCIEcvW48fzMgORks6aE
aFqooOju0PXTuBmQPUHqPJnii5dX1WsB/1hZ+QcmPKgn4QIOpF+DK6NAF7ds8BTPzTUkbd36OMJD
SF34ZcHP+rcl/F7quL3NoG+04YtRhNxF3kb/3joL097qZDqwRhHMojxnUSvFvCaIoZ03fNPBfmbd
IKgOYkTXvJ5sXjFVCGITLNn8ycPU1AYp/cxRF6CvRha07ZqNvSuiNMwNv2QcYcPWEbBlxPGHmF5z
SJM5Zvdgz7D6D4Y8KLlIohxn9zwW2yQwt+dSPgsrLPvLkaJWaEFlHfz8jMNuFSNf4PxE4L9szNUL
A8dDbnW2Gox2aoR/R7ZxJL3kiQHvbga66MjfibpoOpgCAvHRwfUt+30xdJEDCWei83X5z5s/g5D/
yQBAXjbHTDMIpqlh8xI+UpXVqj/J9ERFTJByqKQqRmbymm0D/JsLOsS6C3qcoJjy9F7EA7llZyl8
OQ/ebKU2NQZlRCv7/mFNbTuDLnQyhsJx7bfxHDp34oCD+HInZV1wbfg+bJUEN3//WZta8uq8BFca
1w1VpG6L5x9tzl/+W8ZdbrVvwu+OvT4oQGQgFnvHXrzDi1MpoWevjXvArFfe4scHjkziQXIFwE4p
7QzYRAiu7xD0GCY+y05XFh90w9wB2Y2UFR2FB03K7w2FOaMes+SUMviKCt2o8Zf2sYCgeegHkPXF
PiWJfOdNcc7epkLBByAyaf+LSXdUUHXrpQ1xhmRonS4uhDnhXr3um3/W81UINqJ1VrIgvb/Deamc
XdJVCJ1RlWVxtY0/X6GoZQ+UAx7ChcaNk6wKUH1+JOCO+76W0Dei7638qoJLwoCfnU6TLX0YyPqF
AvCR3VBIuud5SVU4aZgnD8dPWpJcv6pk3ycouJiFAvU1hyDNcFvTcAy0SLzFcyMbdE2FVPXPyM7U
JzEddyLYBexLJbQz+teR8N/YtERjo/li/AxmQpcYWgvn1G6+wbfQMcWRJypCeO8gSuoOsKV2ZgqX
5tONJ4DZxJuhQ72JkMvrJ9zKwIoK3KWP8Oly+4cVKbjlfwxWydtqH2dpGaR11BG30xfCrwOwD0mR
s5PSiZyVTZNfBOs6qaVP9QXI7gOqp7M1P60NULcHqym11/2khVb29bEEtdWeEshvD9K8CrYLeEsP
nD5/ujimghWS+GVRwVkzJZmqhnkpCnf9OtLV0SBl1AbiJqPTqC00kY7QVz20CnP87xyvCK0LtXp1
kjWM7zEw8SwMX0PIkFQi0gsGcL6u1L/RmNXykA/cSzP0HtCdiVjgXnjdeINjDbR2rynGsIallKph
LACCBIiMMwVZTxtnxQ9uuz3sp6FfKN0Y5yPYkweQFw4u1lnmt3UE+Iu7YOj9/zU7NHCihFXtrIh2
t3GZ+xqXh75yJYa7+N9iqQ1fXDnwO0MpVLWHwcXnWN6S4Fwu0RvCypmVUyYv827tyb+/DEY9BY2M
KbMn0Ka5EKpilnLRtUmxM7fexUy2ejkqFGZAOPC6YiEZddROJlQmbr14Mq7bNP6NV9HeFrFwVass
3zY+DJg0CT7vTepQYy2Hv74VX4RoxUTlG+ehmxCE/gg3nxKmWG27GXRje2+mdgheSFxUPe66msQc
iEjiBjOv18bsmmSiebaGvGevSPtYXW8Lk3ihECV/IcYCPPEa2hw948iCGtKMDH9iGJVRN29EIxog
lFBZVVF6c20BEyrw2p0lVjbBdBTFgxZN8OYF/JRB5OQvq3G8gvUZdIx/D1nQgTrvc0Wfvbp1+Uxw
40IRe7BIHefzN2M2w1Ba+RFJ84UVlEyscUdu5MaAsOJwRML8F8C9BB8+w+qTQMD7oJ/eMSLUbWCA
G7OvtjCk5I5JPvhXp816Inj7Mq/tTy3zmgWEaTc1C4zOUrwVbNlNdnL0HRMiX+yGIBAlZ7W7nmTF
314bPgHtvrwkf9haRCuaiect5ePRI1mgYC05poefOpkqhDK+2cQDPRJ4ZEDU5v4SfLDs9i9xO7WI
AR7RBnXjRM7zsJxZ4jkUQeqhaSTN+VR0nMuqW9K9AV0jaRtZfaZX6+029GRdnsR6kcFDg3K363TM
ln59gUZsfjAqB7a3G/ZFhr/Etz2pxV7bXejUrdBTQBFyce5TNyoO1FeSf211HuOc74H6U09eil9I
4VjNeb6uiZiwytDXCMhdIWl4oN7UMEbyKDfCc/qJFXUBXbpHFhSd6Q72GDX5pa7MOKg9CYX14E+k
ddUfQGjJAnK83Y3HBqk2CkhQEEMQwTWsRjK2gvwYrlCi4wdHeMANrPgNWZkDf507+20IBUC6kSAO
5q3oTGM9hSWWbUQCUErUAE8kgHZ7exyshiNmFvmphypZqcbs7muqUYa5Dyi+OX1g+hccpu2DhgvK
FAt8juSrxG49d5T+TJb7ZR/VgKTkkoWFywTHEXMd+ct1y5szjOHjeWpc7egdBBKQZvM4od7R1Pt1
n0cJ7V5PGqi581T+OL8ksDWhsaDcRMQRu78bCaz6IBl6GuN7MRg9BiwL3OaEocgjVAKtFRhZOJaV
3ZnurYHi3sQBeMBzbuC6H3H+F1p5NM3IAbaSRHBrD6gI/Eam5b8MZoGzGNC60He/qW2jIQHeIkTK
fz2HRz//RqVir6wYlJo2g7JgRtMrd6Sq8HyXCMG8bEsTFAB1EqbqcihmPCLmpHdJv2I0Kab/yUVM
kXy1GBTaqmtSS95ta6E4fJIwKPXn3y7VEfYz6hb8jwybiwGXgCbXwuV6he9nxI3E/rsw1c8DpuWO
+NnYoi4dPJ9MV1+oBYqq2XJkjAWj36cvHjLbeUbKy+lDXevU2C3JhzUcGYDnI12R3kdpbVHfEZ7h
EuTd5uAT9MbY8gfj4AEdPY7D5F+TDHWHcuQvm194wUWcx9F9v5ZhGq5NgQ79bQKgu1CvkRdVfWLK
NuCGhID7oeDnFr81iYFoN/2+TXRyoQtAGq3l+UM5WQsyAr9KvXj3mcCjT+g/9jXsiOknjCTMxgdS
Daf2eXmBJ29qfu/lg/sU2LXUx44w9X2hGQkqAz9zYiFqGGl11mRDlqs8EsBIRdY5He5nAC0YYEMm
qlj7d9LP32K+KYuU7/5IWb661TCXwNbpuuRJOhAI0lFIpzTt0tHP0+7nKqwiP5/yqZeNGsnNqtoo
7TbJzFi1lbcwgUZ3pV8KXfk3eZGRJzMvClYYqTBqdH0SmVL+Us9iaLiVh2nAKnvJVpdFJE0kWdYN
aY4T+S7kH9prBRpQzsPSFHHsACug1VnNJoqLPrytcKNmfqgSTKRJ3gqsDn0vX7DM4cV8lzx0CEu2
fxivzdKp4smG3WtXHDDmR/ec4+SXCb4XO1XbUFGP8KjIdbOqiPtkjKYTFlIXnDHYa+zbGk25BJ3b
IFOrxHtDaAz0BNL0KFHq+FsyCmNY+MMQeMKhvtrNsZb+ABq//jpY2ZiJdOSIaF1ON0gmDpOPj3WA
soCePtYEVg9Lymi5BVe2dm73n4CHSiphP/Z2eUrk7T9pW8Y+mGt7xcEwSWfLG/JSQ2I9JeAIRmOx
4lHbMqqr5ZozcXzuH2ans1fQIGzexxz8RjKrBX0g953NwdJ970fKKwhIOBfvXhGBtOYu57orN4Eo
y8gxc1KzTUQCD/RXXtGSigZZnIrVaC9LclpZp1NNhMGd0Q05dsjhMiIK8lZoQkjl52ve751voAWf
gEYTQtD1xrkYAg/pmMHlr5Lvm0kD4naQUxTVXahbuiDt50C2T6t4Tapzt/K10RiLF+Ix5WCUDGdi
vjVOZZLG5xSIbtstVdpn4aOLgh8PwX+ItBxjzAwQT0lal40zjqMVrv+DXvyZ5UeOeKtzmXM3a719
a9xcBk/Vqb8DU0xunsHIwMX8KnDhBCbs40jrUcz2n0laZ5eGW/zGmyUPTvjbMihZlmSui0Kq9Q0I
uK34J8+crA8snXiiLjesLVdpuumelTFKP2WpFYZuVhz7hvQS0l6wESLXYHx6LPhYLHcH/zKmJVjQ
vRg3lmh8ihDtn+WrLpJX84So8ADeYk94GL36MkN1xVcBv5peGZYvKbTeTGldKf4V1lEzLzzk6Hoj
Hj5+hNs3ExWN7pYQA7DVuW+UmRJxfOvuxT2tIer2kr696HjMOx5vIxeRvyhZzyW7kRcI7efo2zKs
wjehgTRIwrG7ooSKU++Vmd0F9EDkEpNjmTbdQ8FxToBWiZNPq7X7DnehLKyPTN/279ig/GkfcO3p
MPdW6eZQnx5fUhjryvWntYvTsW9UK/5HsC0mi28jk8FtFMaz9kw7no3KWzltucSN5sxyiOnqS9a9
Y8y9v2RdseEbAKS6/OkZav3Br6qgpjm3Ryxre5wrY1fPOQMjbYThFcwIFkW8TJqYQ2BSL78Z2UhU
B4k24ROr5xYwSdD7uykKrnDwl3jRYWncVLd/hYZi8Y1zqReVskLRiop8OjTSb0YZYsFfZrsIlbTW
nhcCKcLnxDcyUemD6LAOSd4gw6S6Rs8GBp2ZJCkYwKosiuJG47p8FsNd+i+9vq9MTCnyKCAQ08nd
+r0CeUog26ZkVTZOu4TiTnNF0WLNQaq611d0O/h17CpvDQGPZO1w3njvxtC1WgVOohCTYZwUqWeG
k3xM4TGk5d6Qyuy1dqMpq22j7umlcwCbIE2wYns+EGiBf/k8lWWmVgukR3aPCSvODb3mDuGgfyqg
Ew1q9SPUyG8gkZblNasyeCIMcTnfOo8yNFUJ82+vBeXW1zycYThL0oo+PYb+wjv6Vxv1MIzTJub0
AWNXRp/lfuOYI3bmm+izVlCskT/ex7f1QAGlcTsB2m74NbxhL/xXfdx8sTnlh3xWgOg2lxE0XVq/
jdojV4m/5x7cWyDJulUjlXoK6UoCofENSsya61y/JSKjSakJHsoztMNvkBXDcbAzL/C78vo9NXvU
gtqDngGu/xMliDl7/oe3oHPkIbZ8fKQJwp6pIJoPktiJTYq2p3iIb/5dF6IbS1HIQ/oXUjrWkRUQ
JFey0GuzxQoFOQO7ovGb7lkYGdgMMqqFvKRtoinnJPwmnMrYtcps3X7agTFDf5WNNSMD9gjzG74m
4odmWUzQ2504iD6DwVniSwADryF3M0Bn0oqbyQfkJA0u7tCPraJCosIO6W2c1wZMBrObeVL8ebGj
RO2PSzXlNW45y+HVjDEmUCP8ZNNh4zUvDVqQRm9XJgG5oYpAje+YNJetAkUB5Fo0zSx1aW4o3rb2
GWqG0X02/jCRw3kJ0OxDJ1hOsvfaKrw/wOCLBWeQU11lPP1wav0fk8eIDPla0OjeYJkMBDIpvzEj
l4SdpxMVhJ/ArZvX1FKKAmW3LtXNRA3yAKZgt2lna0xAH5qM2lp40FyvY95Mu09nH175J6BINDqr
cTcQ5gwfLa7mg16Wk+tYJ/D4EVvzgFlghgz0V4UJY94uTfg5wPSrt9jFhHYwxMmzW67VBnxZKwjf
Bu66M61sveqVTxGMdmr2OZaO+lO6gEGkxBoeVnTcNH6GMpIMWqoQKx4PWCw0R9KhpQiUsORc21JQ
aYUcXqP8qoraK8icziWwQgWdtdc7SzZRIQHg8Ple62TngHOt+fGhb2uw/6K/RC9nRsyMlBs5seGX
TvosBnnQZJTNzkSOoVkl7c9IqXprO+CQ8s57GRC8LmOQ2HuSGO4Sjb9M97mPBrkeBbbXE1ASCpAL
LJUIDpAox1oCYnKBKnSAU9cKjyrs1BwtQLrpiJosM8mcWiG6qgXDnye/8EJrYDKqJohKhhbN6cpX
KrgW2WemH7VVOfJfcX4UXyDE8IsQdHU5xbwrOm5BU9j4Jw7xdo3Pxx/4VRU34qG11hsXlxBb7mFI
ehASkh20ehoZD7Fdf5380Nbcs5Mpku8UIFwUzN1PZpZud3w/01tUWWSOmnLo2sH+Yh1T0Xjv0Hz2
G8BpEbi4Nae/FVBJu90I71QolAvcl4BPoA9EXbz1+hFwFlfe36Fmok/Nc0q6BSovw+d9J5DQBhL4
bhLYMMDurgrYYiBy1C6PcVl3dODa8B8RYcYeDpt1zM4U9Y9LXAWoilBycXvD5knNHSdHcf0rNiX9
wxFg9gexIR8wnRoOxpaATycuRdNSHdwa+kVe8/El72b4A2vIj2IBUAPlAQxEbszf6i2moUT8JSpS
EBZmxv0U5VaaZz2bph/THsJiEJY7maWviRyy20YBRaUxR4IpE2c4D6vI/n9ibWeTXXduFiX5g0hY
lo7ZkLcvxifFQjWlBL1alDhMQq7ZwQe0Hmkf8Yg/RKCxXH94lUKwM7u6frYNAgutRFIvQzkuQ7vg
1Ja7p2yja+2CayMOf8WKWSU6e1NpfaSHaBj1mtPZ9v/fpq44gO06MQvUkYuqPDqcNHXaqDPlEsH0
1rFtkGDeNMSwQ9/4ljXG0/HZQgRM5WOGIgET48LJ8jQGCQixzkgc2HFpAhtrU8U61rtE7urU3886
ttjpzEsJXNb9y20vupFSzA90cAdHdbjeXUQqV7iTnmQRPre7gti662kApX54qfeQHWH0+YKl5O8x
HYtkzr5LMHMFGxgUwAQ482fVI3lU3vG4M6YYNJ0ofVpvDItvMXdtwC7S4lyh7ZjiPm9V86/glx9T
i0jnPMhhu/wNXFzIY5BZGxnYXEUpCAALd0cT/eKcyFQwVjzKAPjBf4wyDf7Sm/muU0nmrthMxdio
wT6TdR5wpCwhuddDYSZfQSOS6AryBogAhSzYNZyn1rfcNtC2dEnvVMoJUK8V0SUcy5B1EnhAcXug
2V6FlU1C6oJK2+wSb5BAg/AcvKRaIbYjpNOnSXb4dB5DSVElFUrOYLYfyf2fu5GnqRQfXzveyjKD
3ByxYi0xQ5l2pZlTDYV5VVU6dNRQ8xA+bZscwsVvcMUOkSJPTah9Xnm65rAazelVoqK6t66Q+6RS
7A4oDFTFeGBHq6Q5WYj1Xf7FSmKEWNyF9PmcdieJ2YjkeczpZUmyCgQra/BJjZbzAgOxv0Q86nTi
QV1yK+tSxiZw4nlR677tz5yAp8Rhkthajm24S5remEKGYW4p9OKwmbxEFMC4OdrDvS5RyJN8BcAf
OS3KdzyJkURjY7xmQDXPUvr4oEs408U0Etc0NCYNU5t8TLH9HI3jsCQZEYBsQr6LQe/hzxw/OlnD
RQtLQVzWyKM3UZ7H51oXRgDh9zmE3jOiWwT+4HTaEhuuPz0S03UU2EJWL6NRSroIMYEE2JYBbaIM
0ejm4wXQ+yrPcubSgH5JuWMJbIK1QIgTgSyJduI4tlVkfmYVvW+B6snB8D8Qo82SF6RrjBEMYAOb
/WQTx1o+Qs9vjsAphGnNor/UzhOvN9YoL0ICZE/G8fYwKZzGq+NxWpkiWmvKOGlrm14lBQ+5Yatb
rZ9ZfVRojlyBcZ3uyPnC7WVoiiaUgGB+x78P2Q3OyXxIyCEtpkOrRk9s7yOp3xTb7NK+U/V9iqpq
ZY/5894kyH9QJVvy/5s6ImvQHGAL+LJo2luq1KYlgET66u6tnkCn/rTAt0aSYVBymGnX37hjzHRO
eI1rkmgdU1+5vgCfGFQp480/dIaLiiRmUp9VoidvwJuISjtCShHbyZrYb6j1nsAtP4yBtNwa1LRu
2A7UhEo4ZWGHq611xRQq4f8qR1reIR/675olMUJMquT8Q9cKJhTsMnQroSoNtyG0GAO4mEnvwpjE
NklT5v0IN9oqlkxyeuDf8v7Yfyr2mfw2EmzzEnpwIa8T/gK+nSX+0gMPOtmiPk5TnZkooa4R7s7S
bobb0/nNp0TcKQQDki9lTJz0NJq1L/OVE7swxRXRUqNg3WAyD4H3lDq+7opZKpAHZx030a9xHMbc
yXQMf4fkv6Na84yUWjiY1xomVfNGrioGzYypkS9QSl69x4Q2Eu8TSI0nL0m04mbP9Ec89haulFxl
fPTz9aXI6efQL93pB/YKrrQeHU5K6+iONNvueaKgHc3X0IQpv8OIvksgdgflsyBriwH7LUkZOgrV
pN0IObp4Ut5nzVdO4ZVaBxyEPQrqJQqJWF00ZQKpMBeXM80vLBYxwvU9aLHmMAQk2TQZrOJpL5+y
A5ii3Qpd+7xkLFu+GYoHb8PXGZ7y40yoD2Hr6JXs49yXaHuUDPtmydvJLfvkLqUdvTDGzRoWEKBZ
saCTZxt2GAll6Nz3fxYuYcQtK1AgsqO0ji+ijiXF3/pWB88GR1nJuD1iNPv6sC1wSCtvfbAQ56To
b4IYodTKNDgkWgX75FG180KcPKAtcqQL9PyqgBhEjnDy1Z0HITrcJHHW/QTMyWdMR9k0APlFDUqH
ZMucnW1/tKtxCfAoJFkyLHLFQATyvCH+C7kgY5Qq3EQ4N4v82LEXXBxk6I1osT8T5xLI9uLLMnfH
dU5HDS+wa7PJ0lOyPk6ZdWvHOZARXjAHcKRAHW0fizeHXDgprCIJwCe/bRVjV+nY0i+T4/2YCEi9
Y2RXxTcyADdbye44xdjE+f/fxjp/ppdD0hbgom3pXKJ4S8S1i9HKB0X3LLfETM9h5C16pX5wuZsL
CeJWd7AYbqUr5vu5Vw3zkDf+LE1unAWI53GRxMV68DPSOwg3SMgO74r5UMqoTHZGB0CmbaeJcD5C
yOxh1SkNNui+I3RjkQuu1j1lkNZQ5fcLY/+SB6ll78w2/JKcnqbk+9eja4OJf48x/4sB0QRY+/hv
CgsOBSSCn1jxc5snGqoBmay6PDqCEVngw7D47wEq7Jtrn09GdJ1xW42FWs/bZYcH37/JGI4LoJ6n
DVN5UU78QL1Lx8cKll+b+A08OK2XOFsq01YjsJqdbALKFI1Icx3sp4SY74DSQYr+5Y+rMhtoBXxe
t7O+OoaIIZeJ3vMBtzj91lr178MRbc+215/6Q8nTGvFopnC7N/jjW5P45QfgqTlKPFkNmY1/Tb/5
hrjZc9nELS5l4SbcZcLS3NgwBjMv02Hj8/pa+HJfw3m/YI3AlDY1Sf2Ops5sxkWCB2i3II5sIVfc
yXypNCEmGspCAoE/hDth6C2GFJWr0JezXELa2M2LEOdK4cQeUbriqNC3WrE7CtzA4RCCYDuqwgs6
F4rSPGJYl+WWHEJFYbZSXxEo1LrZFYorDONH68YVks99H1x4H0qkkoWhcajxHKUm6X3mYmTIdlqd
HwNobihQHry1hruQMHSANaLoxOosSRLOT6G2O1uvVzjL0mS8SCXB5Cr2wWqZ+gBpEAUhWlTDArCC
2pDvGvnLGs1wtizRRQ97oKdsZrf6nRBzPAilyJFye0TGjzpps3KNNHO7l1kF9Pyh+1imX67PqLQ7
Cryl3nlaWubbj2Rz1rWFnPri8lPSFCUHFoZ5qkin/K7PFAjCUTpS09AZZlMu1fHPg9GZ2vBsxR+F
DRTGCNaVbugk/BLL1hX28sU5Vg1AhhoF8p/+8EP/lH6h9XUseJ6bo6s8FDFMnYIre5EUjkpurn9y
kNat3o4F8Y9oGWwGLjtauLwqy1Vp3nOzybH2jNhTkxdjyD1WCqSW92BqxLLyGsTXdevqrOG0Yb/7
I8xOMXcaxwvMrB2trkjRdrGFLtOoSEofB2D3pY8b5NPPfb1Dy2/+PNoEy0VgxrBp0RQJdFITnK3p
HNlg703RCP5/ypuik+NbhR+iktxi92jEcTpxpIdHERWCT8Hshs+q3LXLCz76aWfAo36Uhhw54EAQ
ArgXjezdNjT8UKvHj1KjaZSSufbgXeFhzjVPUSAqffSx0RwcPl4xU5VPb6iPQIvNRaG6mIvWbTjX
mfONfTnLawE8ewVjio/vZ+zLzym4KzGeNlqKYSpjGeQEYKaGUYtiYLbwLhs32SrUyP8DYQbq2kTC
09w2opmFZ9zXyXWvXhAOQKgZPrOhbkT+eLhpwKmyASwOQyaT4YupocVSbZgQYyIuNnsVkiJGq8Pa
4id2HUlMeygA/h5rAaOh/DJ+r0dqu/5Plw26oHRc2T3iLf0uRLnADikn+I2xXBWNp71eZUd1Pfxe
dtPQPt5PvmEDZYhOfZpVz/dK8LqqQyGKTrRqnGpXwHHNkinvmM4tE48iQZIKYIHTM2pIfC8u1ItZ
bs+st8E1fKwQ2fwoLO0zCVR7OlghedM4FC5liavyZZ0k1xsOp+e+ktDK2DKwoCJPgZt0VfU39ZGL
ZsA5Ner3ZTf/xDtmOsyUWmIP9XwUby0AXwJ97uHuS3nT0n+RS4mAG7gO7pQdpbK5JNtRDynBd5mL
mquBOKTkjfMHXYs4G8dN28HMk9HTFXu3zBXvT5asNrPucCZesIhxBzM2OGl4zy6hEEVZpwexpFkC
H8BEIf1lIFWwhxONaydMp1TXyCK7HFRrnUK3cMo3ehdtb9UvKAEDpVvEq74iMO6yTVD9VoHPoLGA
dZGjYCojmyCPOBXzpyGV/iFSgCjMHDwtrwE1DPb7kY6OUzb3mCg1bqFrIXv7foPyCbuOa5IvA567
EOgpWnWNREqDxYISmflBreDI+C4BfgCRjMvhtpazZDYydhawHi4v064ms0H6Osb1xK1GanEoIDHS
hBwQ23LmZCSoH4lbJlOpIMPBoZGDtm/4ovG8gBFxD2O5bj/FBSI0iQRlKF16gudfuYjW6qkaml+n
YKtVr4KnjgFdEhotDNjZJ3OyaWu8AFqWKRVnMMs+WXtLlXe4V6mAmbj1z/EAO1lOenFwcCxQqJqm
hKhvWcqi5nuXLaH6Zp5Wy6KQAhCS6vVdbgJ2tjEvHJ2gmaBtCN2Ao6X2tEdRo74nO2YwbaSOBa8G
ixX9ecMTzRkLUh90zpHr4J5fozIrp2vzeff1uzIbip7kksDS/tzK0MA3ZjK7etwseK4ja5/Nj8yS
TYOy60vIWxbUcGPv4aVDD1vrCWbqm40LCRx1wyl3P8H56IgDVTDQ77kZYbXzuIcecCXrmaOcykOV
WkKaYqrIW4UbdjeR9geDI1QLEe1eodwtKTIxMn1Ayp/a6/UIlpKlNYMt+Os8/9M0e4+yeyixF4E8
XR9G4enhC/AI/dBNdq+HG10hqmbWFxzNmq/YF8l/5nyi1Wu3asWKRveYyzQHiJ5l5Q7qkFaFCc+j
C0uJADq4gSQBVbBwl6XVaTQc8O8JMj4ORmKGOmHSBB9Kphto9tWY+Q+A7+TfRePHc4Gaug4Di553
z0MKhsJiNAXlSRBTlovSnXRVKODAw7huYaGRfyWbEKuZs13K1/li2mX+tn06vTbAObDDJj/7x50e
ancBBerAMvQC+u4CgNt67d+7ouyGY/aMQ/WR03j+BxCxpPak7S6RKgy6T8Froa2+AAm/cpwPE/dL
E5Omdhi8L0xoPa5SaaBtCkrB8YPqTFSEOP6WyOF2I+mGjNmApElEZQUMB1o1k3D9GS4l0Rj7rvdt
NXzSkhXbdIxTC7ZyamrhifXUulMcqlQMZ0j88rcEPqNsqToR3PKc52K9IucIkr0Yd3U/c2NlaDFQ
nyeGVapDz4TmT29yoVdc0v+xPtchK8Vkikr5HcH7U8WIxdESJ9FWTuTMfhoS+Ew/eRqQDu123Jjd
+9BH8Gq2RQo7KjnShaaNjlHiA6+gr3WPkOMts2K69src0+zSXtIkWeZgIlRDBABBXVmzM1+IW33N
blyQhnCVVwzuX8p3fHUOfdpbzmmOPy4JwcuW51s4mok1EtTU0C856d9GO+ArdcRmMGPFkvdm0aas
aIp0F9GltBLR6G9aaxzz4or+o7U/wK8w+xKmd2MkVAQHTLbw+y6m3zOXw09nAzJ2TRbXWEOqGU2i
fv3pBuwYKrb/NG5LDrzCjAE5lPvP7Y5c90Id6TaH1Z7i+SISXd+n07QUIl5w4qGHjaKvD5MMhnRL
pucfS3kPxQKcxv+TjoOdyDtwt8wNHM5zZKRSEq14OgvkNCUV7B5FpxPwn8f0pNP38CjMUKeA99yk
l7a2JPgxOY6o3wyeuvlZXLRsGl23Ky8S2EJsGtkm17ecGN3wdBIf4xrZXxIFoAHw+aEq8Ta+rbjb
8mucwMrveSGOwsW4Ol+t8TNmH1lNxWWpaXSgm5bDY2dO9CFMHvIYDBVDmLYrIh7nxSATjfWuIUwq
dZ+/d75HF1hhWjLp3n4BDFV/MvppHAm9SsZoJOxm6FTXp/lmMXp7BjpqgV8ptQK9cB/olkRkeegT
YyAGSdVZua/s6UkLSV5E4VAeO9H95L58Ax2fFWWCoC8bFyVeCurfKq7DOgD4/fIRbZNRtm8iZO5V
7h1TfhPrmxvNhRx9BHQbnrd6+plGJiCfQ3bhR+0phJF1Yxb6wDq67Hp34hfOiRfl3b3D6+38Ua2/
dquwRjBUzcvi99RTP6Pe7DpOdCOA5QOu1ihfE/ttvfOHCEenU57q0vPvGGbv9ifusbVoLzadA5rF
92J/xfX/T+iOy/tniUHpNtWkxQoCyDbZ2uqeCRT02OaMTfLcQsWVP346Q6HvIDUtKdmU0OSCwnZm
yKYmdP8uCsw8ENB2jg/wPragz5bsRX5SqIHyZ/94ptwe1Rk7JxPzwpGz2nweQxzcv/MT5g/necMj
NdfQSYo7/8NgzNqcJEUrGRtJsHNP2fgjbufxy+WtD/HGfcD2jtX+AvVrKCBTQe9hN+3dcqCJ0CB+
tqojFjGF1jeHIOrotBUC1L3/QtMaAygj06lhkeFWIrkdhiXnukv8caauq3rKFHIeNQFEF/8PdMTe
p6M08U6J869uYJCaV8ua2ZqnnOZTLQSYGhz7t2u8ZGSTpIABbZYowE22xWC4Ng4YNJM1vIe6GBxv
KN/QiiC8KZQWlFuWelV1EZrLXAcnxFje6NKJ3I/lg/82IzMViqRnBJAkccQC7bT6o6pEyA8p2qmq
51ZSTQ+rEheOhKm8plduvoVYkq8lOML9/tK/Y2u0BOW1EiOig7MIIdlqJDKcrq5EubsMzOaeeZf7
tUMChQJkDlv19rtUc1woojpmMM6gIfVLmuJsAbKQr7BT8zVmoU5o1xPK+TCPBsfrvydIjBKxvbbY
bxG6aaLf5iwXMkzAxVNsg+K1aehDg+jjBgW3dw2goAgZTsejENJNukIsLWQatkBpdK8kYlrE7SWv
ivyCpMRugPACgS/WhjpNjS5zyeANoFNMnM/wR0wdvMro1yOd3HGvZR4OWrqJ2TtuKqm7oNtUhmol
qoB4zyNZGOk1tGd/OtTjXE3iW887/ki3Si8nsieGI8sNfilP2fu+Z6ljhGKjN7E4ZHWEfHOcQct3
R1KJz0bltp69Yl5VQEdtA4R6cWriUmyR3IHHfgwE+AMhHXcdNXNVhB3u3D2X5TREjsdVrpegymI+
HmWha3WROs8gxiPV7yC62DX5Wp3xfP2e2mUcH55MrtDVi651hBGgIM2yAkrAerlrsp8XSlxpt5xa
m+NJrcQ9wL9QixTSrkJtbuTGCJkMMikmpVKZXSd23i39lb+d9X9dKZ6kc4p865vCJ1JczXMcwVrz
0DcuvgFeeAndGLHhpWxbRIAh2ISe07XWGhloJQFp5C2PCmAn7wjGMqAbwUKpusGEWfD33tnraAlY
T63TJrf8I92PKs48EyO9Tkyu3Wd6iA/GK/nM8S0FbkME1k5NDKGb7xtFttGYg0KgSNgLuYupHDHt
UA87GxHxe1u+20qwbX2Jh5iEL/k91sGi45ZujzwlfG5qnTaFEGkjV935Xpvx7/luOUM+qMEvJ4He
ma57jQYkbxvrJblbeNBFgVU6YIT14mbLokxB0P5KCLHGWDX1R25JqnK2fEMW6M5hKAzDkBByICzK
nkUCSfHrffOULUNzMit+yO+etNmd03/OSPbCK94zLf5vmLdo51fmJOOQ3Ep+3k2zIUbrfKr6QZiY
B1mZkT8SsLgJ7x1DtdGHs7lQ6pr+Ko67GzxULbRFTYiTrsfniIiun47N5RQh2E67/cxwT/ouH3hD
2xNMfmMPGjwO2JeBbGmmvezgYzBaxwJ/+97YaA8pRuGOlLoM7ma1tprNFLwzLtVMi80fnUEHYxIn
dq+29eUXf/uD9gcH/Hxm5L6BCosvXh4IhD5tkhyjwE3sOdrHFskmNbddfGQJumpV6tJ5sEP0FAkC
bMfL01saLljff2gwq7bfiZXzJgGU6ZI2iBm5lfew5G6G4Bdo3usS6OQdtfjmSHS29ySJpRRwH9cq
GQ2iUt2Tcx6O7Ulx4HStfUp0gWTcRnO3/8B3qHkpnL+gzACxysxzWx+l7b6dJVjPFvAIYqjADUTT
k0G8oiaFFTESe9as4vkpFj8emTY6ZrT4ndPO6QO9ZtSku9p2sY92T5GmZw1BX9iTJDTsm+yOrJsT
hOUSrJ8uzFeTCqnlW1QUa+fI3R4gZ4uIMtFXLOq34ohL2SGF80/wHFKHv28Hlknp1dBPPfVBp82T
aBMT73XKB+xUQCMF6LSxyIuiFLbr+Tfe6GJug4T6mxwH5U6t2c/tqFk3JsKhAzjvVQRxhbFNOSfG
gfW7fPdFASe9WmA6HnspBDWVSxbj/KUEtXW44OyEZqrCBCOchN/AIAQjrKNt60qi9OnQEhuXZCr4
ZXlH165FWXGSr3ynb+xa+p+gT3RdNXVgFp1ZshRtdMagN5uLOqRFTxtS0x0kIZyC/rw3CsLZ/z09
liaXAxeDR4VpT6zEs8EDSrmw8lgAkkC/EuDKO24tP/rtSz4wVgp1R5HubjIFQwZ7Hxea5eqwtJIa
Y7CYH84L2gZ7VIi2Np9s9pbBhLKnDszG56FJ8t/DqyBux1ALTyjq3OH3U1CvoWto1phA2NXnmrl1
RVe3/rUdOghvZ1cY5I3HTv2pLA3VCj4+ewAjdQPdhq2czMgs2oEobBUM9MKRWvMdkRS7uA9/M3qO
sQCX5d2RtJNcemmvy5LoYTxl6LXAhKcLibvvST7Z6MEKOI8ZTr7O4bK1KjOGIcmApyE/iTkS65jS
DVnoBR2p69v7eQUcRPXJRJdS8tkw7toBIGLixPUbEg2QPxQ5poCe3uP7Cpci8oKk1NAcjFkQkQrG
EodWqOz1Al3tNGbqJVQwR47Of84hqEnbQ6ji4Knfg1rVQ1KNgWout7dFjr8lAhFTq5FBY15Wb/Jq
jdiLU0jNNYggVUEHrY2QKBDNGTCE6eZVKYDDY8gnPNgh0xqsgDYyUOuxmzlrQ+o49D+L8A/BkAPh
UBn+/DBh/gkeukme16VRe/XRHDsqdHm6boP88YmMYFDuhQWIosT7RzUt7TaFrQuVB9PJ1lEAFa+6
typGtXx7DofjisnPHFpKXbE0nYB1FT+UThX8LGx4OjtsKEysA3Uox7J5xIZb3JyNS1cx+MCqCPW+
NOgMiXxzRZeJC+8Eb/RFGeMdIm2h9chfxCM5GVy5lyopfKBtPCHi6yNhU9cqST2sACugaj2/PHjS
3lCoIsEzKSZ5K2YHQiF9PrKRKEBCPgWztZUO4l9hvye2+XAHsKJsqajQgTHlcZpryPjudX+KTD1J
hwugK+km0+Y5E0qI1SxJrC4q+Fao0ceemFWSgHf4TEeZk4ci5vDwN+CP4hPin09gLkM2xHoRpwJw
3TD7864cfpJxkZbnGh3CuS6Y7g+kK6Z7gzALN4u4ZjBV59fhxh99XQpM6/lNcCE+UJLCA8rxm2wI
zHQrUBBWWaw94fEP4SAbfGI5YiJ3cnPAqKXWD1PCMULMGajfG0Qwq7d1yygzGojacW1TSgS/mDNT
QcaqA8NyxgVkC+NdB0q+WK5xJB+Lf7APic2bf+9+Iaweum1iLOJnwChWz1g9lIkATUxUXHAvVOrK
GMT5awgWAH92xtLAXWmQoY81Wn225+1e4aVUBFf5TTKVvvhBQnFHwQLbjfnUqovt0zk5Ga0eqFfW
UA75Np6yWAH6386iIo7scNWklRSXsvsu2Her/B2hLrnneG0MH6Cj5p82ifIexh3F6Hs+OO/7CQdG
N/Ff96Bg14vPaBIzT+P/5CYtwX3I5jgXrI+XaYKd72RRdXWQUEmVjdpttuceuEXR27052Vj4WPRR
4rvTmbvpy79TDA9sQwkgDGQfxbuHFZdQft+P8yrljp7fFCHJfX6U4VdPOvWF2I6FpEbvzfIs+gDq
eFtHe76bCmr8kU9A8ONkLDH2KGkSOrKO16NXy8sagvqhKyaTtb87IhAPw0TmbhaMGsC+R00t4JR1
vlTk7jbEPfhG+pHNs4S+e8gk78IIyUMX09zEdlMiQBnxPtwlwkrrZcbHAkaxuWz8z1JDYF2wV7Dz
CnzfNLltGJU/tPo5CwSqqgbPPu/ZhBNYuX7328+3g1HSe58Vh5noVy8Ip+hcQpOg9jDvG83uw8nv
nyu9RxtFbdFrr86rer5Lrh3n7rmB3iM40gQhuQAZLg3lM+xooMsU3iGgM9lNbNDq6Ne+0r3J2+sd
ir9QJlVDfNzNpmxs66JGKnY3NE80TadJQ8LhBbX+slohkoZlqgttt/OhhaosYC0Oxq4tNvps9S8v
tu/G0XRRObjzNaNUMDlmaBznTsLJHiVGyuX0GUX6NHxP5GYDwo8L7hXkbxcySzMviXu6aGGjW2UY
40pBS/4wz+KlvRn5cODZS4Ypjb6OThHv12Aa3cUN+BFx+sSU1UhinCwC1mpKTA2Qh2DTg2CuWppA
t43wH6olh+6f1Y9AKIjdXf335eAdZmk6/XboJVA0c0iKkH68KF50HQkUxL4Ji1E4lttFfEnM4Bt8
M12/3sb0Dkz25Q9SNljbyMh1YSr6UP9bKQxmqNkkS5mOedwmMsKVpdYrYFhPosXLwPoHHC3dNu2V
n56l9KuF+UfnRdu6phjsb1APgTsyLn0TgDPFaAQbb1kdhEHFKUDzuYs0oTmaNGXHGHSg30rnY3m6
IZFaWf8e5e6pQv1TP8D919Qob4J0gENtwV1TKKTbXAm4zFDg2ebA6xq708wI2bpWuyFP6MEHY+BI
wauoAjvzsZvqUIHgJXtEXZibmhgC1uSWjcSev6JhDX8Jaqb46EEVxUm+ayYJdEqeILEMjQt5fkUK
dLUzi92G2dKNiIZX4JYnbv37E7CWsjYaCrRQLUW5VWThfwGkw88bK9Bcx+kdVKcHlxpcqRPQxrLK
SPfk1jrGASnqfXfnHn+Ogtf1O9c7AgWYMbEsOOZKo/5IvlPT403aufsaXQG0NDEDDQjVanRmAxN4
XBtysfTNGdXD9fulQlgzHk3AWD6DEbauaRoCss2FPdyrsdwRNbn3J2M6nWnyu3oyJaLSP+NHZewq
z8P5P0MNOYi5f/e9aWUsoutPp8U5gicSo+CX/h4uUKgpd8eOGVaF03Jj47JV9sORl6JPyY0BnjqP
gHEKUB/anvdR1NdGXb27aAoruMhy0C4mm11vfi2bvItwaMHN2ESpug4NoK3zJJsAGBE4oE74OFS6
zCapgSl20bFFYIyaoBUFC3m2ggyiKgQEYL6aBe3YFtk+9SuF+hx60K31x0Y35kGFj+6ji91xfD3B
jeOjwICUz4F5P7rDFsCpeU10FJtf7TpfJBchxu7Q5QAASiQIKlGlzWNwWWx31D/d/l/B3AEtu3DL
phddV7q+E0x1uJ8dKIEPZR9Qs7+QPnhF3tQmZpfiUH9YgzsF1CxG32kOHirJdSCMx8OPQyUml/JP
VlBdC9hFeiSRJOdnaegqjrhBTje7DreBeaZ2qw00pu9VzrsyT80aANHqbij0jy5J4Fsu3+QM1/cg
5anvSgTkG/UmPcboo1AQ32ZLV9X5IPP1HelnxagpG07fpA+neXVDW/XkmazgvGxoz0xtrMcVhs5D
qKsfq5BgMWsyfdQtdk8vsZQCInE8/lcbUt8UHXcRlme5P2IQ9/vvgkMBn5J/r/mJmvcJY9p296lF
zklOfrEhVaqNinwA/eBXMuhJ1QMJOJsKJTRujG5OMyyToya7jIxNQs5ozmXrEk2bHdcB9QP70ykm
P+ZDeDZ7mGDYBDo9abt5OZ6+NV5bjoNoVLBEpjrZnB0KcBR1/6i1/DNhiWOxjZDcUfKUIP5EOkKv
uY+1g2n1COl2Q6GRIFDF4tMr1CdPfFfWGR47G3EShO5vQJ402iBjNWdLD/O7zE4dzGlZPCyH38yH
Uwi5hsQ+RFP21QxPYM+MebvBymW7KWZ/E3CZY+TB3blVaK8hpWAteXqg1tYfqVwfwR5MMsm1W0Aa
gbrhRjgri0mGio2eky+ZJtuqDkc5O1OOxmvFLYkpKta4x2D5OUfI0It/ShTOg3GD1z6qcS60mnqH
ypRH0sec5gMkKn2ctsHwp1CWBkXipdcUDgHFm8EKPKFLV54Lg7LkIn2rjyuGNcKEyffgDseQhxZ3
L/A196g4leuXJcI8WfhqfRBjBk6z/Z3srurYhBCzLAMnkLzRumKV6ZEV68V/pqXuktlPNukkhDdZ
gihSKG1baavyKBXFjdJ7nOYfr4ZDOp/jSSlD6DfM2mbf7ITcTRmmZRiNKXCN5qfyEDTUsfoaOysN
HZ8ZBfNa28jQmHeL3OwyX+9rh9rxCc/geMNvRsYtegQz39SNOJooRjlgztOvaZD/3/61WEXTKlQR
6J1XnOLV9kWm2N/IUjPWxiwUJZJyvchqza7oczYfYjX+Lo2bzAYECbyz0GttTJvztf3Fao6CMp0P
HhunNoHLT3Vtmf8xL9mZLFGMRSySRjMw9VyOntC22Wl7OgpKoY4Xvt7GyEohG240U1PSbNJYd5Da
L22xDuh9RUGT3604iQbYYIp4CJsonwhbWqc/ojEdr25RDFoWKn275IzSQHsE1d7Hls/Ex6DyHjZo
qLLaz9FqpenYNA4G/T7lFfo3YPygaoQ7np8gFMpv/6u/dQQ0fGzjrcQwA+JbcfSUelnU84jVKds1
fT2hZyDx8hbv3etnwzzQWc1XzRzhfgCREidULCXHX5MkSB+CImJCoDByiGQl6uo20WI03bUSLF9B
a6iq7ECXN2Gbi+O+QwUBiz1ne545p0GeiTFtuWtetwbu7hXdaFGPBz0BCdm0jp/Kfl1lfRbON5pg
NlN1UFcAIQE5OvJeqyS9lOX0YaeeijhuMAgj9KuNFO17HKG/eF/PbOrmUVuVLn1bd3ap2KFzZQvE
MR7oKGoNdlTSXs5gJXm+aOA4F25cS5ZEWNjTzfXQoCCXNgI8tibMbRlyEcfykZ/c2on1DtIiYafV
ixB+ZQc2a3UrcUBi05RiXSVPQm41//tObMLAkenmymjZW2nw/NjFrM5mKutoiNAv6EwfuPkcGnS3
CmT+EmDPr5DgyEQU3g9M/Qdhv/YySmgSAeDoPJZ0YkE0LhCwmzqqWewE+j9PViY5+t7SvgoXxTnY
BabHb+oIezLdua3TV+DnevIe9yK1pv2rMZ6s7MLqSyxRknBL0x+s18nbcqDnLyq8ENUveJD4RitN
BnD1WChx5RN08lMg6bzSSFyHzOkXZ6LxH+xRrrIKtmhjGT1bCNADlIzzyoCFKRKf0+ZZymova+OW
iQltjYj+EpsFtEYNlJJZ9BppnzQpzjkf5mN0co8KIHTgdYXgSECzuwx9suN3vbDYm2wzQp9UJ85z
vmHBHjqzxKdAFj6Ai0cOn6f2u3SP3dC61DoWg6smHDNqMgfYp3dBVYBcI63NiDt89fjLjmwVyo+i
yOB+4bChCt2Hnl3NknTAVy7+RctqTGjgn/95nYzqGX1V0k65dsw9FIMSqKSsxtEnkmRfoFF3aTRc
gULmcyYYWg4xuiWHEYAujGn+6WhJc6fE6HSDvJRXHPGBy6HIS3sB6mGNqz8Uh/kl5ma7Z3OZ6GyJ
X7SQFQLhuYBSP/ygCMuPzdwiZUemMvegMJVbgmlpl9vQIXmDwXG0VXbUxWrAMIjPpRfz95B+hsI7
kmYMxLAyxR0PkLNr/0IujnQJoRJo1jlX7M5awsTCIrGomVb5MwHhtkcp4JmC7MAwQg2OecvMD/hS
B+rCRvA5qDHw+JAnyO9u09iXEbh9sV6E6EhfUZHQB9kMd90+RmiNIksBimhV/dqePW1PvP5pFbX1
27egCnmfUJ03juJxB1yJeh33Cq4u1FiHwR2/AOPZJxu9xQAJCfXBBsOHMzEetGwIkorI1ZFfCj8u
vv9V7XtuEYvjgnWpfydrBXn4BeenAJ0nnFGO8+86ixFutynn8h4mAp1r/maNBMx9DP6WSnw4ip22
ZrxgsKe2JgsUFAbyt/HwsCbn+tGum/tNt1yLlIMtPuquTDL1xWsrrwMvE4Y9d13mReey2E6OdZCh
G/6iTgapr7TfFfaXVn8SrPftCXZp0diuuB1pXDIMKzjn8y6FSeT4hMBj+zHbHBIdLqQ4ZZG6LqiI
YR7MCSI95pW3yZ+Y6ayPQB/tXqgMtokCFYxOXWR0B9Jwjz1Wgqv3dMIe/oRO2fpL5JPckxjw1fI/
ombeRByt7gizEKYWpoLtQGgqndyM9TSM1CuMtb6XnT27eUUiQo7+piVsyplN0NyvEjPRzHnJrVRw
oYW+9XngWQ7Oo4kFA7RFbOs9fQj4daL737kDxpEC1Zg7C81var0LH4OwanCL2twcLZrF1aYu2u7z
qBdCsR/Lr5a4ENNDcY6gJY3Dc8A37FypPNb0SXwpub2pCHEj2nOZ3Jq0XU/vGVvYe6xDCHrkn0Gv
p9Q0XO96B3to2mPANRIGleBrs27AkdwF2ZxqsZnAG9Fh9UCrs0R03GddI9RJK15TA0FoCFLvkkQT
UbUxfXzdBS4ivvDtbyiRG5wKrpuHPz7FwBxSRocT+1h44eCjSUpPZsPWgCtuUG45s6YZUSQzSa5x
4Uz/qcBjIKVHs2qE+kzeJJE+FfOvv+MP1JpclZUYqH4iaphWOuRotgWsbQYMR/qnm+E+w1mkc1rs
VpAzACRDhqE17pvxNulNtcXWNDNYtZM6vW3yCSchyak/yEkW2ShHnj/EPq/jW2D8tZ5qvyWhsQx9
7cIwa1HlTB83VZchASKmD7+17VlTHzJs4hCAygITu6CJxQicrj+5FTB3/TnQfpTJcb49J1XZhbXj
+khrLxvL0h68a5JYglS5SQtJaLRhQlrVG3ruiSw3hFd0nP+r+l1d/7tkSEutbnDOAOpvYzcTqyIf
Gtq7l166j4rfaq9be+pCER4rWzZncdba3O1QZSxoXRvDFkQ5dNK2jyqBO0j5ta0iLDzDXvn85Ehb
Lg8UJ6EdCBL+azMNJZLAmDOzIlJhrRuNs7BMSIIlQaKNTUBKlscVRez2pYz3hDWo00JsC8jByk1l
/Jq9o6qTwz36pIlfoFUfTtwzFO6a6Grzt6kC8dcs45vvRJoOdKRPmNi6EE5asvwz9e2i1x1k3PM0
pnIrKJtYUnroIRkl+Q0xi48L3/HiSkiTAuiAgae/hSmazswHOvFqyFxZNJfAB2UDvk+CISthMx54
JueZxnvCSNKojwiQrIlD/KLji5SmJNNfmYOznYKgYiGnA1kQLbW1nLQVNp/5S1FZcctaMZmJh2x+
cr/tlqJdHr703fRlwwmJtU3okdD5LRwjMP/EeufnSRYdWBDeX9Oqu+as2k/caINBuWUrO/+gUjwA
EmMqsfMgov0Z7uvg5/L38QXAHNEi0wvOBhQXi7g9k78leN0tJmyE2aEntY2lysuIW0xXN4drD3E5
AfHBL6F/LbwelNpisNFJ8RvdwXpVdyutyOb9dmm3yf53rFVZ+426mwpzFTUwcBBcC76NHCrDHaz+
sb5/J/NSj8IDd/FOh8chZ2LlmTlMzuu2pwPQbzgrt/ewG6zwmjYnV5l1SDlI3jvKoQt7uhnKd4RL
LiEm9wiHDd3IPhK0mz+fPYtc6rsvAMiP3Epm3EdBwlEsqUrjltLDqMlf1VOjdSdL7oRLyAfX3e+f
BjgEp1l2+SXY2R07MF99S0Lukl5Aa47eXimrx5Rj2zC5MWrdjicSgNTfLMlcuLCekTaPff9PFOAG
QVKdyuMxYasSnTBLhE7VsptPCYdw4rtbe5qrlaACFEE29bP3dHInyixR3r3ZqymY+WOyKJIU4UMF
TBmTY5nFyGpet3e0N1yCkKjah8Ff/uHrfGcHZcJLWMeyWq61u4mBx1agYIl2tYL1nvcTvqf5XaZT
uMlOGngaOSbSQ6dukx/rPwq2VlUaJ7KWC0s/RjXgul2Yb5bnG14wtSDZ6FOJr/LIucMEV6EFY5s5
lP1tOOqSDp0K+XyiTsTyfZs3rLEp0MAZpCyUkCBjsQQIz+7+RfTGhKTNl59O71BYRSud3RHKtU0I
pBiSPQXdPJWQUqZExjLAEi9cy4DlwxwosHFGgr3KWnfmXaP9A12CxP6cgPX5YVYB7DQqhCNo84+a
TrhqrOQa7XDrX2ksOkoK5Hxk4dW9pzJuzMGZixaNSRSOwSHxcSUriMi/15DH0er4v7lLXcy+sN0i
ZiOohH5mGQZ1uddw+RT6S0li6Qv7rEb1hJt4jajvN2JnmXjSHQ4fxuk6VDtYuyNU+CFvJGuUz8vf
SwZGWML/2nfh93z/kYFjqgNYBTy+4pzbs/2bqlEo7nw3weV1uRHNv4uxXnbPim5Tqpg8Q5m3vlzg
g7g1Eyk6wZo/Ywl9YkHvIop76Rxdiw4l2ngzxOw/xBZE+UKUQhanO7O79azx/otnUmtn621z0Dtj
0iJClZDvXz7P50OFtj3fy0Av3kisTDzJ4KEzD6S2ytZguu6ySMXtBa7NlbbNQsaA9f19UG3Iww8S
luQkh5LyxE6lDMM+lmFpQPlucZ4J9coMclFOlBeGj9wkBTVmzOYR63jW2LG0XJed0ya6QFfyy2i0
JLVN8nlHV2Y3kNH3Z+zJ2wxYHckGXi3e0/BYTLZivDk/DazhHOQjufTXN7hqwdbs1uFzn3Fgt7hR
6GlCQ788ZDb6Cuv02UMwtKb53leEVZdYgyUMqKrlS/dc7ULRpbGjOsQV37z7wc0red7Y3EBpsUbi
U+X+ZY+Dw6QmSVtj4YtvRewLt5Hh5kIAzvUrOuFil2wBq8EomTz3AxuUq/w816g54arWObtNmTix
ABv1GMipIA548PeDLUULfTRtyi406XEyXdoW8Idxi8gtRSIPRTCBJFscQqviASl1FH1heiaYA1cU
dCD7qikydz4J11xzJ4+y92ylNWdirGktGb8mlzrgkyTxzvWG7UasDGN31cVYsdk9QXQt1fz4iWVC
Du34oYyYSQMMGdGJwovIxrzC7aAqeWNJi8J547PKOic3lyZKfqWiodIE/ZEmcKjyAhzeHk9BBzE3
lRFtUDMOmH/XOZ2htKfSfNe9BYkvuwg+RVjj+DA9I+wjf8rFUK8PKsGoEVwx5XV6i5G9vRqIDYG/
rqeBbzYSCb79Z8G7hF15gAogcmpWwrPhta9AjOrJd91/bprZb9lBg5zPL/4XJiiKMbjSVEOWE8Q7
9Xf+5pSp0gTTSXl0N4CXOiqg38e9jiI8nFKCX4KYDwHEJbAohsK+KLsYiptWW+xC2aasfTuNcPfj
5e0Lc7kxGwaHTdj28PACeGuEtWoGd10ond5L8tZZo19pYxPGTLMwZEmmP4WhIZVJLQihOCQ5/Xdp
Wp9QyJeDGz4O47TQ+EpeMNjLbUDoZzZZFTVYmsHHpdXnpgbBBQ101JLlX1dG9hiBV8E56ONDIxBP
Rjz3QfqWJLv0VVdYjdaTcWVZHq2r0r/GXEIQ8MJdEXHr2G6psoIZK6t9Fyisvdt9MRPdy89JdgCO
b/JhBwiR0sHNGtCorUZR4xZQTOR1gvbDujX1ibmxkVOB/t/1ecvi08DNLq+t+r9ltHScicmnOiJe
nsHFvZXuitS0GXvYJO+mqX6ywlSKO0NHIE355M5P0cO5qnEDjWb8uXRf6IyCQzGz6LNyb+upglz6
n38LnKa5/h32g165YF/dvl29Bg7DGOhKHNmgCdFhTvXyQxbARMFtdaP09/MFloEPZIwzWo0FcTJb
MIlWWqleyXJMpH2xhw6MCk0tc/nbergS4BaCtzTL5ZCXSffSMmdmy98AvYy5VXy1PDGYZ1CveAXA
0xVjbBV5zKYr2cpPbW4lvIenUdAWLTquz1VdsFFgyvtTZKL+thyOk1p6+ZJPgJZdVxep2NilDfR8
E6IfbdYgcXbhhAnjXZ88BxXkrA0RQjmL5cy+6Iur/Rz4NNELPIS9g23uyfDU0AiQAr7u0bSOxYUb
0ddnd9ZGU+XCGgbpGVd8JAkxzibP6TnPPnJBlf8Eqg5Kkenh4FxdHtCrB57nFuR3Dli5gBoB+bMc
+gKkYXLDpzsg2dQvL+iq1iPjMBgBT4ykBEv8qnLnmf9bGESvnT9UYRhowAr7yv0JOfrSoJm8ctlg
ri9ow6Z397MQLWxuQvP4Yh2dZ8fSaL+Bom6vhWe/1a5Nhn0DgsKUjRbXqJZ34N0i64KD9BcA6oqm
t5QuENHO+TX8C94kbuMcmOsrQ7rVzYpCOeBC687MLGN+6Fj0s8Af/8yesA+Au408oqlWZjuQJlyd
BiIpyygjOsf3y180k0wx1wu4hbUd3N4o/Rz88gtWhfWMZlSn2G904ONTCD9jle7sYEL/4BKdcsxN
HQOhbVxoIG0oQu+Q2hU06JMLZWa7xGma/IGqNBeiPQtwtWhQZdyLQcydbRp/oE+GGzUMrVA4/j2U
VgkiSujH7WZm+pIO1AtdF2UqXSsICD+N+qG2HYNCsbEWBRjLIvJ7D64BSlBTaZ1Fwa1RrC0DjWf+
Rr2vCVGd5Uu5RtX8WzHaerujaGcFfB8XaS3jll1R2bZqeJ0iGYKR7RAch+N9IcQ30EUd38vEbO9O
wzRm/kZLdIE34T5tr4FsbOAq+V9NqhECYQ3/PK7CQOzsMJDUcRd42oumtgx0mbhPy2rPD5ECLLQf
avi+uai1vz/wbFESFK2eSPjawaCvV9tSF2IY2vbCVCHDCXMO2bye4KuxeeYq1kVjUmXgWnC4tSL5
g7VFwfc+qV3s8YtBrcL9S9LTKIcoduLuwwKvXB05l/osCvZE/ee2YPZ+YORkhmWlfSNcAsdeQija
98ndm4hbwQ13A72JuA3QW3yd7Ombx2uj7dukcAbk9rz9PWhTGlHDRsl/OkUovSEt1ADeb3APY6J0
AIXkMHVpTgUZPGO3lcfqF6pgxVd3PnkrZrPHM87FFH/p9MwwXisQTd+hjeNxG8DO6l4yC6bDIHD3
bSUH/Vare8g88BhOcP0WZ44p1Ofj27pHV4qiNFaPyimQRSnrxGLNwtXfiYORrTqmJm+FwcPN3vfH
uWM5jsfFiY4f4Kn1A5SObqHlGo7Ui9j6gYTRYHOSg+PTNUBv2FL7CFk36Zby6KReMQoifdtmkzPd
UdEfqMdyBUJs3A4P9lXRAjSExys0hdkjaqgtJWYzIEjqc8LJi5ocMUWY6tjQAT9MgZqrzsEsOIp+
X1AWJjNOQIXeHvu0irovPMj1V0XzKRxp7pD5EhMTH70dVrZfi35CZry5VVsMTmZNxH1jvJPJrvX+
utMjt1Z7fql7bskGy7c30NXqYKKmtQZeTHc4XL0WhZm7qu9n4GGFS0VMcvAiF4kFOKJCwFLJdI8J
/PMsCHg59+vMqTl3LOMjIEyy4hmN16rdvXpIlADfGGLEeIRQPrRxgWZ5k/gEegqCOQKYRYGfz7OQ
GgxF6UZftgy7b/m0WGL48vOwtlru/vC0+GGbnebtzG8D4Fa95Epb8oehyf/6/WDfjo8UWFQV4Tpf
FVGQkppfDkPkdX/qLBScebbvhswd5jFHPBZh+J3NQWrvfwQ/DGsKqHJ6TGpiG2r2b7j+8TIBsLIL
tLeaBJ0K3Y3Sjr7aPpajTCEo3fzXq3WAtI3lus+o/Z77bl0DzE3JhpMqL0+COcJkGKgbnmcn7akh
YcmkqO8R3mZsJm5hm/cxy+fFJS/7Y3kaR+ZpImdtvfpx+AOcQD5pIyu/rLCA6wxbjsWDlS4LqZKU
wHi+7yudOewC/iIFHosHwE6WL6Ug1LnwVzsStJGPjMt/YJhh30320MsCE1yEVOzqnCUdKvCWm+iA
tY0W/SeYqChR2wZR9tQX0C4kANiCgtkHxfzVxQJrBndnrWrP8Dh5zHAoivcKYCga9iPGtD6ehsVC
EyPPRw+Ripum2rommEWzMDCsmRPc2ZI1JUgECmQIth1JUakPBPXj0GqXAepdHDfo+2Ku/mwQks1G
Klbxc/asoL8Suj0n/82bKsJFDkU9juqwfFL42ZYvwPzeCSzy60Kszat5SYFeW6n65+JeL0rvO4zZ
Fg7CDVQrJalW5SRXedZrvtfu9NEyFDVKfRnHfCn1W/2EOWW+OZPc5u4OMBpOUlIkJ5cTSWPmEwq/
iMu9peNWigVMvfxdivljfW5lLaX9pkjTIJTWpalaSNl/B2RudurnEpzsv7IV+A8YixVEGwyt1wNG
Gsd6fvHFDpUStrbubSa7T+LSAIlffsFW+EhjXQZPgLYpolDiSqzzD525zQt7D2Z7N5knHK9Pllbb
rJZns33OlqwtuZs64YkUX3OJ7FaQ/zQuv3u4bfTp0/gZmBelNT1DKr6vsboCa8PA7LjzAn0PK0DU
uGtdj/Gpfb4i7mEa7miBi81FA33oLQgJpDiadH0o+y4ZQMkQyEbntvt6nOBfr0NQNt7JZr13KHaH
Y2PtG6Fs3ylwq3+bDPJvC1EKcPz+/IZKSvV7by7do0IFGUMh5gq96aGxa0kjCEETdhnMVSTC+6Ax
81xy8/K1NS0Fy6BY3budxqT+1xaC3lLQQwMDOZEz8OmNgjVqycrBeDeXx6k21ZLMzdp072JrDdKv
x4RsJUomSuFZhwmaHmBme+jfMp0ExvKw+Ea7QL+MgC+Ud3K/e9fI3nYEf/mpyJi5Pe74qDhMdh5l
zXMwhNFgHvHYtFuiQfdX09OLvIrcOePtxm8+N68vikasw1stFiTe/Vn+dQUc5Raf2c0V+ewb9bo9
kFqOEk/y2zSR6QaUeMS5b2XydaWZutJtUaLe+dAJ67RqolTiCwILT3I1/3xPEnnXLNG7BajFPER+
fmafG1iAeFMZO4cUv4g2iLWxHk62MvGhXN0bvY9nDAKSWqGlwAJa/lkZlwj+jIWn9Rqk+5VHE/eU
+551VjGXBjNaU8oRmZ2MoPAx6eUD9laVQVQMr9eogLe0pT6qz55wr13Ohxy+h3Cyc3UGHciSF+sG
GYNKH9o/4BZDo5Fb5/Ujw1pJBP+Q7oBNzHMHABPU0cUGK9Y96IR2k2eIXA0omgY2i/GSjGi5cbTg
nQReGDFh71muI3+tgiwyGuzWB0bDmdtSKuTj4EaCmq0hD2y6H46yuu7MJ0+MXs0YftySFvrxMI45
F20+VTzVUPLkxxk1bpPLHXQWRRmUlM5IO1A5W1MSLEjyhocLMvrgUAJwjWHVkgPG1Lth9CnQ0K79
Oqm19mgFsC+JlhRcalWqNII+FDRf+zezLfHENA+tuEKT5Lai/+oP3iwLXsy/WLAzOECASsvHJF06
L7Lrxw9iWCupVhy67pXys16nyseYRlc8i6NDREjDaRcWxE5+DouYURmVWMXK6m0TYAiJAsPEs9ra
hqfe6IRRpFWJeiqfdQlYxGV6Mb4heLuUIC1GVIGRsJLIh5vqSKlgZLbn4fBhmeWwSZPEPXV2uCn7
363jVlJctPLtPZJ3A3P3QAnQtImsC3uIN7DP1wT5ylmzQj6sseHKDq9OiJYExi+r2JBACZ8tVPkZ
QVa9dJwSjVCCKmb/OelcRAfjghC6Kzg2O4pVE36BPBlvB0l0tM+R8YSd5ti3zHL73taSNuN5yXBB
wmXLgMXrAOFlioegvQ0OV1IV1oRQ14EhBEQhhB3/rsod/oABai1F4w49krfq1Cq3ZmZ/qMQ6EEQS
FzEBM5Yw0SoJVZOdGUGg1lZV9mJ3UoenTcGT3R7SIR3g6Y2kFybMcZQRtzRr3Ph7VwhOt0MUVSEn
xp5aBPHZLISP0EyUkdehzgqb+1UBduK3M4/9AfLtL/cGPHeell+a4higzJ6Da7IewjCiIrMNfY8o
qgfwMh33PmHBMwRHuzrdwVVe/Kt9J6/ThaNUuFyznTHjqF/3e5OmAXdpFPDWws+ZKeuqyJspzAEJ
MeoJYvGttOhja8+NjbszscQR4xVom+MEULWE1i4/YcOUy6oxVGd3ZFU/0vtw7f3vshvOv8r46NUn
jwb8YhgveoapauvCChLi1xAwflA+dIUzVwRGJnx+jH+nJF91PJW1yXNOW1LdJ4IQkx+3cPK1V8fN
dhKRGla2P2bHIm3TbjK9kiyLuBm0bKJw5cHua6+wc4buHn6Be1bQ/KRrtaDM/xdJB6heaS2lzvhC
yvGxng5SR8ldsPE7UcKO9UJ1nu9A5y1/L6b7ulQVJU/l7DntInhNB6dM2ou/zPuzTc+uSYCODVir
SbKdbafJUbduA3ZgIOZwEnYuf0Abn9aGywZJ+P7Jbk2vDuXDDZCNN1Qf2yDopLXrdVKsXKk1mgy6
oOvhywwd3CFGiAKfYsy3yuECR+JxhUvDHRSC/7x9p5UP5RUvj2Rfsfe7ESglf5RlK/beSmgjsxlv
r5gL2eSa2VUI01hXrD2Ctz8JASDtQYM83nMMHixxcZJCThBdKMLJlNRNfujXnruQSaPDQJSEr2d0
ErHloQ==
`protect end_protected
