Package p1_pack is
Type sh_reg_sel is (no_op,load,shift);
end p1_pack;
